module krnl_tsp_rtl_int #(
    parameter integer  C_S_AXI_CONTROL_DATA_WIDTH = 32,
    parameter integer  C_S_AXI_CONTROL_ADDR_WIDTH = 10,
    parameter integer  C_M_AXI_GMEM_ID_WIDTH = 1,
    parameter integer  C_M_AXI_GMEM_ADDR_WIDTH = 64,
    parameter integer  C_M_AXI_GMEM_DATA_WIDTH = 64
)
(
    // System signals
    input  wire  ap_clk,
    input  wire  ap_rst_n,

    // AXI4 master interface 
    output                                  m00_axi_gmem_AWVALID,
    input                                   m00_axi_gmem_AWREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m00_axi_gmem_AWADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m00_axi_gmem_AWID,
    output  [7:0]                           m00_axi_gmem_AWLEN,
    output  [2:0]                           m00_axi_gmem_AWSIZE,
    output  [1:0]                           m00_axi_gmem_AWBURST,
    output  [1:0]                           m00_axi_gmem_AWLOCK,
    output  [3:0]                           m00_axi_gmem_AWCACHE,
    output  [2:0]                           m00_axi_gmem_AWPROT,
    output  [3:0]                           m00_axi_gmem_AWQOS,
    output  [3:0]                           m00_axi_gmem_AWREGION,
    output                                  m00_axi_gmem_WVALID,
    input                                   m00_axi_gmem_WREADY,
    output  [C_M_AXI_GMEM_DATA_WIDTH-1:0]   m00_axi_gmem_WDATA,
    output  [C_M_AXI_GMEM_DATA_WIDTH/8-1:0] m00_axi_gmem_WSTRB,
    output                                  m00_axi_gmem_WLAST,
    output                                  m00_axi_gmem_ARVALID,
    input                                   m00_axi_gmem_ARREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m00_axi_gmem_ARADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH-1:0]     m00_axi_gmem_ARID,
    output  [7:0]                           m00_axi_gmem_ARLEN,
    output  [2:0]                           m00_axi_gmem_ARSIZE,
    output  [1:0]                           m00_axi_gmem_ARBURST,
    output  [1:0]                           m00_axi_gmem_ARLOCK,
    output  [3:0]                           m00_axi_gmem_ARCACHE,
    output  [2:0]                           m00_axi_gmem_ARPROT,
    output  [3:0]                           m00_axi_gmem_ARQOS,
    output  [3:0]                           m00_axi_gmem_ARREGION,
    input                                   m00_axi_gmem_RVALID,
    output                                  m00_axi_gmem_RREADY,
    input   [C_M_AXI_GMEM_DATA_WIDTH - 1:0] m00_axi_gmem_RDATA,
    input                                   m00_axi_gmem_RLAST,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m00_axi_gmem_RID,
    input   [1:0]                           m00_axi_gmem_RRESP,
    input                                   m00_axi_gmem_BVALID,
    output                                  m00_axi_gmem_BREADY,
    input   [1:0]                           m00_axi_gmem_BRESP,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m00_axi_gmem_BID,

    // AXI4 master interface 
    output                                  m01_axi_gmem_AWVALID,
    input                                   m01_axi_gmem_AWREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m01_axi_gmem_AWADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m01_axi_gmem_AWID,
    output  [7:0]                           m01_axi_gmem_AWLEN,
    output  [2:0]                           m01_axi_gmem_AWSIZE,
    output  [1:0]                           m01_axi_gmem_AWBURST,
    output  [1:0]                           m01_axi_gmem_AWLOCK,
    output  [3:0]                           m01_axi_gmem_AWCACHE,
    output  [2:0]                           m01_axi_gmem_AWPROT,
    output  [3:0]                           m01_axi_gmem_AWQOS,
    output  [3:0]                           m01_axi_gmem_AWREGION,
    output                                  m01_axi_gmem_WVALID,
    input                                   m01_axi_gmem_WREADY,
    output  [C_M_AXI_GMEM_DATA_WIDTH-1:0]   m01_axi_gmem_WDATA,
    output  [C_M_AXI_GMEM_DATA_WIDTH/8-1:0] m01_axi_gmem_WSTRB,
    output                                  m01_axi_gmem_WLAST,
    output                                  m01_axi_gmem_ARVALID,
    input                                   m01_axi_gmem_ARREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m01_axi_gmem_ARADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH-1:0]     m01_axi_gmem_ARID,
    output  [7:0]                           m01_axi_gmem_ARLEN,
    output  [2:0]                           m01_axi_gmem_ARSIZE,
    output  [1:0]                           m01_axi_gmem_ARBURST,
    output  [1:0]                           m01_axi_gmem_ARLOCK,
    output  [3:0]                           m01_axi_gmem_ARCACHE,
    output  [2:0]                           m01_axi_gmem_ARPROT,
    output  [3:0]                           m01_axi_gmem_ARQOS,
    output  [3:0]                           m01_axi_gmem_ARREGION,
    input                                   m01_axi_gmem_RVALID,
    output                                  m01_axi_gmem_RREADY,
    input   [C_M_AXI_GMEM_DATA_WIDTH - 1:0] m01_axi_gmem_RDATA,
    input                                   m01_axi_gmem_RLAST,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m01_axi_gmem_RID,
    input   [1:0]                           m01_axi_gmem_RRESP,
    input                                   m01_axi_gmem_BVALID,
    output                                  m01_axi_gmem_BREADY,
    input   [1:0]                           m01_axi_gmem_BRESP,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m01_axi_gmem_BID,

    // AXI4 master interface 
    output                                  m02_axi_gmem_AWVALID,
    input                                   m02_axi_gmem_AWREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m02_axi_gmem_AWADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m02_axi_gmem_AWID,
    output  [7:0]                           m02_axi_gmem_AWLEN,
    output  [2:0]                           m02_axi_gmem_AWSIZE,
    output  [1:0]                           m02_axi_gmem_AWBURST,
    output  [1:0]                           m02_axi_gmem_AWLOCK,
    output  [3:0]                           m02_axi_gmem_AWCACHE,
    output  [2:0]                           m02_axi_gmem_AWPROT,
    output  [3:0]                           m02_axi_gmem_AWQOS,
    output  [3:0]                           m02_axi_gmem_AWREGION,
    output                                  m02_axi_gmem_WVALID,
    input                                   m02_axi_gmem_WREADY,
    output  [C_M_AXI_GMEM_DATA_WIDTH-1:0]   m02_axi_gmem_WDATA,
    output  [C_M_AXI_GMEM_DATA_WIDTH/8-1:0] m02_axi_gmem_WSTRB,
    output                                  m02_axi_gmem_WLAST,
    output                                  m02_axi_gmem_ARVALID,
    input                                   m02_axi_gmem_ARREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m02_axi_gmem_ARADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH-1:0]     m02_axi_gmem_ARID,
    output  [7:0]                           m02_axi_gmem_ARLEN,
    output  [2:0]                           m02_axi_gmem_ARSIZE,
    output  [1:0]                           m02_axi_gmem_ARBURST,
    output  [1:0]                           m02_axi_gmem_ARLOCK,
    output  [3:0]                           m02_axi_gmem_ARCACHE,
    output  [2:0]                           m02_axi_gmem_ARPROT,
    output  [3:0]                           m02_axi_gmem_ARQOS,
    output  [3:0]                           m02_axi_gmem_ARREGION,
    input                                   m02_axi_gmem_RVALID,
    output                                  m02_axi_gmem_RREADY,
    input   [C_M_AXI_GMEM_DATA_WIDTH - 1:0] m02_axi_gmem_RDATA,
    input                                   m02_axi_gmem_RLAST,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m02_axi_gmem_RID,
    input   [1:0]                           m02_axi_gmem_RRESP,
    input                                   m02_axi_gmem_BVALID,
    output                                  m02_axi_gmem_BREADY,
    input   [1:0]                           m02_axi_gmem_BRESP,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m02_axi_gmem_BID,

    // AXI4 master interface 
    output                                  m03_axi_gmem_AWVALID,
    input                                   m03_axi_gmem_AWREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m03_axi_gmem_AWADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m03_axi_gmem_AWID,
    output  [7:0]                           m03_axi_gmem_AWLEN,
    output  [2:0]                           m03_axi_gmem_AWSIZE,
    output  [1:0]                           m03_axi_gmem_AWBURST,
    output  [1:0]                           m03_axi_gmem_AWLOCK,
    output  [3:0]                           m03_axi_gmem_AWCACHE,
    output  [2:0]                           m03_axi_gmem_AWPROT,
    output  [3:0]                           m03_axi_gmem_AWQOS,
    output  [3:0]                           m03_axi_gmem_AWREGION,
    output                                  m03_axi_gmem_WVALID,
    input                                   m03_axi_gmem_WREADY,
    output  [C_M_AXI_GMEM_DATA_WIDTH-1:0]   m03_axi_gmem_WDATA,
    output  [C_M_AXI_GMEM_DATA_WIDTH/8-1:0] m03_axi_gmem_WSTRB,
    output                                  m03_axi_gmem_WLAST,
    output                                  m03_axi_gmem_ARVALID,
    input                                   m03_axi_gmem_ARREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m03_axi_gmem_ARADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH-1:0]     m03_axi_gmem_ARID,
    output  [7:0]                           m03_axi_gmem_ARLEN,
    output  [2:0]                           m03_axi_gmem_ARSIZE,
    output  [1:0]                           m03_axi_gmem_ARBURST,
    output  [1:0]                           m03_axi_gmem_ARLOCK,
    output  [3:0]                           m03_axi_gmem_ARCACHE,
    output  [2:0]                           m03_axi_gmem_ARPROT,
    output  [3:0]                           m03_axi_gmem_ARQOS,
    output  [3:0]                           m03_axi_gmem_ARREGION,
    input                                   m03_axi_gmem_RVALID,
    output                                  m03_axi_gmem_RREADY,
    input   [C_M_AXI_GMEM_DATA_WIDTH - 1:0] m03_axi_gmem_RDATA,
    input                                   m03_axi_gmem_RLAST,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m03_axi_gmem_RID,
    input   [1:0]                           m03_axi_gmem_RRESP,
    input                                   m03_axi_gmem_BVALID,
    output                                  m03_axi_gmem_BREADY,
    input   [1:0]                           m03_axi_gmem_BRESP,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m03_axi_gmem_BID,

    // AXI4 master interface 
    output                                  m04_axi_gmem_AWVALID,
    input                                   m04_axi_gmem_AWREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m04_axi_gmem_AWADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m04_axi_gmem_AWID,
    output  [7:0]                           m04_axi_gmem_AWLEN,
    output  [2:0]                           m04_axi_gmem_AWSIZE,
    output  [1:0]                           m04_axi_gmem_AWBURST,
    output  [1:0]                           m04_axi_gmem_AWLOCK,
    output  [3:0]                           m04_axi_gmem_AWCACHE,
    output  [2:0]                           m04_axi_gmem_AWPROT,
    output  [3:0]                           m04_axi_gmem_AWQOS,
    output  [3:0]                           m04_axi_gmem_AWREGION,
    output                                  m04_axi_gmem_WVALID,
    input                                   m04_axi_gmem_WREADY,
    output  [C_M_AXI_GMEM_DATA_WIDTH-1:0]   m04_axi_gmem_WDATA,
    output  [C_M_AXI_GMEM_DATA_WIDTH/8-1:0] m04_axi_gmem_WSTRB,
    output                                  m04_axi_gmem_WLAST,
    output                                  m04_axi_gmem_ARVALID,
    input                                   m04_axi_gmem_ARREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m04_axi_gmem_ARADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH-1:0]     m04_axi_gmem_ARID,
    output  [7:0]                           m04_axi_gmem_ARLEN,
    output  [2:0]                           m04_axi_gmem_ARSIZE,
    output  [1:0]                           m04_axi_gmem_ARBURST,
    output  [1:0]                           m04_axi_gmem_ARLOCK,
    output  [3:0]                           m04_axi_gmem_ARCACHE,
    output  [2:0]                           m04_axi_gmem_ARPROT,
    output  [3:0]                           m04_axi_gmem_ARQOS,
    output  [3:0]                           m04_axi_gmem_ARREGION,
    input                                   m04_axi_gmem_RVALID,
    output                                  m04_axi_gmem_RREADY,
    input   [C_M_AXI_GMEM_DATA_WIDTH - 1:0] m04_axi_gmem_RDATA,
    input                                   m04_axi_gmem_RLAST,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m04_axi_gmem_RID,
    input   [1:0]                           m04_axi_gmem_RRESP,
    input                                   m04_axi_gmem_BVALID,
    output                                  m04_axi_gmem_BREADY,
    input   [1:0]                           m04_axi_gmem_BRESP,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m04_axi_gmem_BID,

    // AXI4 master interface 
    output                                  m05_axi_gmem_AWVALID,
    input                                   m05_axi_gmem_AWREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m05_axi_gmem_AWADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m05_axi_gmem_AWID,
    output  [7:0]                           m05_axi_gmem_AWLEN,
    output  [2:0]                           m05_axi_gmem_AWSIZE,
    output  [1:0]                           m05_axi_gmem_AWBURST,
    output  [1:0]                           m05_axi_gmem_AWLOCK,
    output  [3:0]                           m05_axi_gmem_AWCACHE,
    output  [2:0]                           m05_axi_gmem_AWPROT,
    output  [3:0]                           m05_axi_gmem_AWQOS,
    output  [3:0]                           m05_axi_gmem_AWREGION,
    output                                  m05_axi_gmem_WVALID,
    input                                   m05_axi_gmem_WREADY,
    output  [C_M_AXI_GMEM_DATA_WIDTH-1:0]   m05_axi_gmem_WDATA,
    output  [C_M_AXI_GMEM_DATA_WIDTH/8-1:0] m05_axi_gmem_WSTRB,
    output                                  m05_axi_gmem_WLAST,
    output                                  m05_axi_gmem_ARVALID,
    input                                   m05_axi_gmem_ARREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m05_axi_gmem_ARADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH-1:0]     m05_axi_gmem_ARID,
    output  [7:0]                           m05_axi_gmem_ARLEN,
    output  [2:0]                           m05_axi_gmem_ARSIZE,
    output  [1:0]                           m05_axi_gmem_ARBURST,
    output  [1:0]                           m05_axi_gmem_ARLOCK,
    output  [3:0]                           m05_axi_gmem_ARCACHE,
    output  [2:0]                           m05_axi_gmem_ARPROT,
    output  [3:0]                           m05_axi_gmem_ARQOS,
    output  [3:0]                           m05_axi_gmem_ARREGION,
    input                                   m05_axi_gmem_RVALID,
    output                                  m05_axi_gmem_RREADY,
    input   [C_M_AXI_GMEM_DATA_WIDTH - 1:0] m05_axi_gmem_RDATA,
    input                                   m05_axi_gmem_RLAST,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m05_axi_gmem_RID,
    input   [1:0]                           m05_axi_gmem_RRESP,
    input                                   m05_axi_gmem_BVALID,
    output                                  m05_axi_gmem_BREADY,
    input   [1:0]                           m05_axi_gmem_BRESP,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m05_axi_gmem_BID,

    // AXI4 master interface 
    output                                  m06_axi_gmem_AWVALID,
    input                                   m06_axi_gmem_AWREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m06_axi_gmem_AWADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m06_axi_gmem_AWID,
    output  [7:0]                           m06_axi_gmem_AWLEN,
    output  [2:0]                           m06_axi_gmem_AWSIZE,
    output  [1:0]                           m06_axi_gmem_AWBURST,
    output  [1:0]                           m06_axi_gmem_AWLOCK,
    output  [3:0]                           m06_axi_gmem_AWCACHE,
    output  [2:0]                           m06_axi_gmem_AWPROT,
    output  [3:0]                           m06_axi_gmem_AWQOS,
    output  [3:0]                           m06_axi_gmem_AWREGION,
    output                                  m06_axi_gmem_WVALID,
    input                                   m06_axi_gmem_WREADY,
    output  [C_M_AXI_GMEM_DATA_WIDTH-1:0]   m06_axi_gmem_WDATA,
    output  [C_M_AXI_GMEM_DATA_WIDTH/8-1:0] m06_axi_gmem_WSTRB,
    output                                  m06_axi_gmem_WLAST,
    output                                  m06_axi_gmem_ARVALID,
    input                                   m06_axi_gmem_ARREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m06_axi_gmem_ARADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH-1:0]     m06_axi_gmem_ARID,
    output  [7:0]                           m06_axi_gmem_ARLEN,
    output  [2:0]                           m06_axi_gmem_ARSIZE,
    output  [1:0]                           m06_axi_gmem_ARBURST,
    output  [1:0]                           m06_axi_gmem_ARLOCK,
    output  [3:0]                           m06_axi_gmem_ARCACHE,
    output  [2:0]                           m06_axi_gmem_ARPROT,
    output  [3:0]                           m06_axi_gmem_ARQOS,
    output  [3:0]                           m06_axi_gmem_ARREGION,
    input                                   m06_axi_gmem_RVALID,
    output                                  m06_axi_gmem_RREADY,
    input   [C_M_AXI_GMEM_DATA_WIDTH - 1:0] m06_axi_gmem_RDATA,
    input                                   m06_axi_gmem_RLAST,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m06_axi_gmem_RID,
    input   [1:0]                           m06_axi_gmem_RRESP,
    input                                   m06_axi_gmem_BVALID,
    output                                  m06_axi_gmem_BREADY,
    input   [1:0]                           m06_axi_gmem_BRESP,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m06_axi_gmem_BID,

    // AXI4 master interface 
    output                                  m07_axi_gmem_AWVALID,
    input                                   m07_axi_gmem_AWREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m07_axi_gmem_AWADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m07_axi_gmem_AWID,
    output  [7:0]                           m07_axi_gmem_AWLEN,
    output  [2:0]                           m07_axi_gmem_AWSIZE,
    output  [1:0]                           m07_axi_gmem_AWBURST,
    output  [1:0]                           m07_axi_gmem_AWLOCK,
    output  [3:0]                           m07_axi_gmem_AWCACHE,
    output  [2:0]                           m07_axi_gmem_AWPROT,
    output  [3:0]                           m07_axi_gmem_AWQOS,
    output  [3:0]                           m07_axi_gmem_AWREGION,
    output                                  m07_axi_gmem_WVALID,
    input                                   m07_axi_gmem_WREADY,
    output  [C_M_AXI_GMEM_DATA_WIDTH-1:0]   m07_axi_gmem_WDATA,
    output  [C_M_AXI_GMEM_DATA_WIDTH/8-1:0] m07_axi_gmem_WSTRB,
    output                                  m07_axi_gmem_WLAST,
    output                                  m07_axi_gmem_ARVALID,
    input                                   m07_axi_gmem_ARREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m07_axi_gmem_ARADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH-1:0]     m07_axi_gmem_ARID,
    output  [7:0]                           m07_axi_gmem_ARLEN,
    output  [2:0]                           m07_axi_gmem_ARSIZE,
    output  [1:0]                           m07_axi_gmem_ARBURST,
    output  [1:0]                           m07_axi_gmem_ARLOCK,
    output  [3:0]                           m07_axi_gmem_ARCACHE,
    output  [2:0]                           m07_axi_gmem_ARPROT,
    output  [3:0]                           m07_axi_gmem_ARQOS,
    output  [3:0]                           m07_axi_gmem_ARREGION,
    input                                   m07_axi_gmem_RVALID,
    output                                  m07_axi_gmem_RREADY,
    input   [C_M_AXI_GMEM_DATA_WIDTH - 1:0] m07_axi_gmem_RDATA,
    input                                   m07_axi_gmem_RLAST,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m07_axi_gmem_RID,
    input   [1:0]                           m07_axi_gmem_RRESP,
    input                                   m07_axi_gmem_BVALID,
    output                                  m07_axi_gmem_BREADY,
    input   [1:0]                           m07_axi_gmem_BRESP,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m07_axi_gmem_BID,

    // AXI4 master interface 
    output                                  m08_axi_gmem_AWVALID,
    input                                   m08_axi_gmem_AWREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m08_axi_gmem_AWADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m08_axi_gmem_AWID,
    output  [7:0]                           m08_axi_gmem_AWLEN,
    output  [2:0]                           m08_axi_gmem_AWSIZE,
    output  [1:0]                           m08_axi_gmem_AWBURST,
    output  [1:0]                           m08_axi_gmem_AWLOCK,
    output  [3:0]                           m08_axi_gmem_AWCACHE,
    output  [2:0]                           m08_axi_gmem_AWPROT,
    output  [3:0]                           m08_axi_gmem_AWQOS,
    output  [3:0]                           m08_axi_gmem_AWREGION,
    output                                  m08_axi_gmem_WVALID,
    input                                   m08_axi_gmem_WREADY,
    output  [C_M_AXI_GMEM_DATA_WIDTH-1:0]   m08_axi_gmem_WDATA,
    output  [C_M_AXI_GMEM_DATA_WIDTH/8-1:0] m08_axi_gmem_WSTRB,
    output                                  m08_axi_gmem_WLAST,
    output                                  m08_axi_gmem_ARVALID,
    input                                   m08_axi_gmem_ARREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m08_axi_gmem_ARADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH-1:0]     m08_axi_gmem_ARID,
    output  [7:0]                           m08_axi_gmem_ARLEN,
    output  [2:0]                           m08_axi_gmem_ARSIZE,
    output  [1:0]                           m08_axi_gmem_ARBURST,
    output  [1:0]                           m08_axi_gmem_ARLOCK,
    output  [3:0]                           m08_axi_gmem_ARCACHE,
    output  [2:0]                           m08_axi_gmem_ARPROT,
    output  [3:0]                           m08_axi_gmem_ARQOS,
    output  [3:0]                           m08_axi_gmem_ARREGION,
    input                                   m08_axi_gmem_RVALID,
    output                                  m08_axi_gmem_RREADY,
    input   [C_M_AXI_GMEM_DATA_WIDTH - 1:0] m08_axi_gmem_RDATA,
    input                                   m08_axi_gmem_RLAST,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m08_axi_gmem_RID,
    input   [1:0]                           m08_axi_gmem_RRESP,
    input                                   m08_axi_gmem_BVALID,
    output                                  m08_axi_gmem_BREADY,
    input   [1:0]                           m08_axi_gmem_BRESP,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m08_axi_gmem_BID,

    // AXI4 master interface 
    output                                  m09_axi_gmem_AWVALID,
    input                                   m09_axi_gmem_AWREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m09_axi_gmem_AWADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m09_axi_gmem_AWID,
    output  [7:0]                           m09_axi_gmem_AWLEN,
    output  [2:0]                           m09_axi_gmem_AWSIZE,
    output  [1:0]                           m09_axi_gmem_AWBURST,
    output  [1:0]                           m09_axi_gmem_AWLOCK,
    output  [3:0]                           m09_axi_gmem_AWCACHE,
    output  [2:0]                           m09_axi_gmem_AWPROT,
    output  [3:0]                           m09_axi_gmem_AWQOS,
    output  [3:0]                           m09_axi_gmem_AWREGION,
    output                                  m09_axi_gmem_WVALID,
    input                                   m09_axi_gmem_WREADY,
    output  [C_M_AXI_GMEM_DATA_WIDTH-1:0]   m09_axi_gmem_WDATA,
    output  [C_M_AXI_GMEM_DATA_WIDTH/8-1:0] m09_axi_gmem_WSTRB,
    output                                  m09_axi_gmem_WLAST,
    output                                  m09_axi_gmem_ARVALID,
    input                                   m09_axi_gmem_ARREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m09_axi_gmem_ARADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH-1:0]     m09_axi_gmem_ARID,
    output  [7:0]                           m09_axi_gmem_ARLEN,
    output  [2:0]                           m09_axi_gmem_ARSIZE,
    output  [1:0]                           m09_axi_gmem_ARBURST,
    output  [1:0]                           m09_axi_gmem_ARLOCK,
    output  [3:0]                           m09_axi_gmem_ARCACHE,
    output  [2:0]                           m09_axi_gmem_ARPROT,
    output  [3:0]                           m09_axi_gmem_ARQOS,
    output  [3:0]                           m09_axi_gmem_ARREGION,
    input                                   m09_axi_gmem_RVALID,
    output                                  m09_axi_gmem_RREADY,
    input   [C_M_AXI_GMEM_DATA_WIDTH - 1:0] m09_axi_gmem_RDATA,
    input                                   m09_axi_gmem_RLAST,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m09_axi_gmem_RID,
    input   [1:0]                           m09_axi_gmem_RRESP,
    input                                   m09_axi_gmem_BVALID,
    output                                  m09_axi_gmem_BREADY,
    input   [1:0]                           m09_axi_gmem_BRESP,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m09_axi_gmem_BID,

    // AXI4 master interface 
    output                                  m10_axi_gmem_AWVALID,
    input                                   m10_axi_gmem_AWREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m10_axi_gmem_AWADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m10_axi_gmem_AWID,
    output  [7:0]                           m10_axi_gmem_AWLEN,
    output  [2:0]                           m10_axi_gmem_AWSIZE,
    output  [1:0]                           m10_axi_gmem_AWBURST,
    output  [1:0]                           m10_axi_gmem_AWLOCK,
    output  [3:0]                           m10_axi_gmem_AWCACHE,
    output  [2:0]                           m10_axi_gmem_AWPROT,
    output  [3:0]                           m10_axi_gmem_AWQOS,
    output  [3:0]                           m10_axi_gmem_AWREGION,
    output                                  m10_axi_gmem_WVALID,
    input                                   m10_axi_gmem_WREADY,
    output  [C_M_AXI_GMEM_DATA_WIDTH-1:0]   m10_axi_gmem_WDATA,
    output  [C_M_AXI_GMEM_DATA_WIDTH/8-1:0] m10_axi_gmem_WSTRB,
    output                                  m10_axi_gmem_WLAST,
    output                                  m10_axi_gmem_ARVALID,
    input                                   m10_axi_gmem_ARREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m10_axi_gmem_ARADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH-1:0]     m10_axi_gmem_ARID,
    output  [7:0]                           m10_axi_gmem_ARLEN,
    output  [2:0]                           m10_axi_gmem_ARSIZE,
    output  [1:0]                           m10_axi_gmem_ARBURST,
    output  [1:0]                           m10_axi_gmem_ARLOCK,
    output  [3:0]                           m10_axi_gmem_ARCACHE,
    output  [2:0]                           m10_axi_gmem_ARPROT,
    output  [3:0]                           m10_axi_gmem_ARQOS,
    output  [3:0]                           m10_axi_gmem_ARREGION,
    input                                   m10_axi_gmem_RVALID,
    output                                  m10_axi_gmem_RREADY,
    input   [C_M_AXI_GMEM_DATA_WIDTH - 1:0] m10_axi_gmem_RDATA,
    input                                   m10_axi_gmem_RLAST,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m10_axi_gmem_RID,
    input   [1:0]                           m10_axi_gmem_RRESP,
    input                                   m10_axi_gmem_BVALID,
    output                                  m10_axi_gmem_BREADY,
    input   [1:0]                           m10_axi_gmem_BRESP,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m10_axi_gmem_BID,

    // AXI4 master interface 
    output                                  m11_axi_gmem_AWVALID,
    input                                   m11_axi_gmem_AWREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m11_axi_gmem_AWADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m11_axi_gmem_AWID,
    output  [7:0]                           m11_axi_gmem_AWLEN,
    output  [2:0]                           m11_axi_gmem_AWSIZE,
    output  [1:0]                           m11_axi_gmem_AWBURST,
    output  [1:0]                           m11_axi_gmem_AWLOCK,
    output  [3:0]                           m11_axi_gmem_AWCACHE,
    output  [2:0]                           m11_axi_gmem_AWPROT,
    output  [3:0]                           m11_axi_gmem_AWQOS,
    output  [3:0]                           m11_axi_gmem_AWREGION,
    output                                  m11_axi_gmem_WVALID,
    input                                   m11_axi_gmem_WREADY,
    output  [C_M_AXI_GMEM_DATA_WIDTH-1:0]   m11_axi_gmem_WDATA,
    output  [C_M_AXI_GMEM_DATA_WIDTH/8-1:0] m11_axi_gmem_WSTRB,
    output                                  m11_axi_gmem_WLAST,
    output                                  m11_axi_gmem_ARVALID,
    input                                   m11_axi_gmem_ARREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m11_axi_gmem_ARADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH-1:0]     m11_axi_gmem_ARID,
    output  [7:0]                           m11_axi_gmem_ARLEN,
    output  [2:0]                           m11_axi_gmem_ARSIZE,
    output  [1:0]                           m11_axi_gmem_ARBURST,
    output  [1:0]                           m11_axi_gmem_ARLOCK,
    output  [3:0]                           m11_axi_gmem_ARCACHE,
    output  [2:0]                           m11_axi_gmem_ARPROT,
    output  [3:0]                           m11_axi_gmem_ARQOS,
    output  [3:0]                           m11_axi_gmem_ARREGION,
    input                                   m11_axi_gmem_RVALID,
    output                                  m11_axi_gmem_RREADY,
    input   [C_M_AXI_GMEM_DATA_WIDTH - 1:0] m11_axi_gmem_RDATA,
    input                                   m11_axi_gmem_RLAST,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m11_axi_gmem_RID,
    input   [1:0]                           m11_axi_gmem_RRESP,
    input                                   m11_axi_gmem_BVALID,
    output                                  m11_axi_gmem_BREADY,
    input   [1:0]                           m11_axi_gmem_BRESP,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m11_axi_gmem_BID,

    // AXI4 master interface 
    output                                  m12_axi_gmem_AWVALID,
    input                                   m12_axi_gmem_AWREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m12_axi_gmem_AWADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m12_axi_gmem_AWID,
    output  [7:0]                           m12_axi_gmem_AWLEN,
    output  [2:0]                           m12_axi_gmem_AWSIZE,
    output  [1:0]                           m12_axi_gmem_AWBURST,
    output  [1:0]                           m12_axi_gmem_AWLOCK,
    output  [3:0]                           m12_axi_gmem_AWCACHE,
    output  [2:0]                           m12_axi_gmem_AWPROT,
    output  [3:0]                           m12_axi_gmem_AWQOS,
    output  [3:0]                           m12_axi_gmem_AWREGION,
    output                                  m12_axi_gmem_WVALID,
    input                                   m12_axi_gmem_WREADY,
    output  [C_M_AXI_GMEM_DATA_WIDTH-1:0]   m12_axi_gmem_WDATA,
    output  [C_M_AXI_GMEM_DATA_WIDTH/8-1:0] m12_axi_gmem_WSTRB,
    output                                  m12_axi_gmem_WLAST,
    output                                  m12_axi_gmem_ARVALID,
    input                                   m12_axi_gmem_ARREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m12_axi_gmem_ARADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH-1:0]     m12_axi_gmem_ARID,
    output  [7:0]                           m12_axi_gmem_ARLEN,
    output  [2:0]                           m12_axi_gmem_ARSIZE,
    output  [1:0]                           m12_axi_gmem_ARBURST,
    output  [1:0]                           m12_axi_gmem_ARLOCK,
    output  [3:0]                           m12_axi_gmem_ARCACHE,
    output  [2:0]                           m12_axi_gmem_ARPROT,
    output  [3:0]                           m12_axi_gmem_ARQOS,
    output  [3:0]                           m12_axi_gmem_ARREGION,
    input                                   m12_axi_gmem_RVALID,
    output                                  m12_axi_gmem_RREADY,
    input   [C_M_AXI_GMEM_DATA_WIDTH - 1:0] m12_axi_gmem_RDATA,
    input                                   m12_axi_gmem_RLAST,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m12_axi_gmem_RID,
    input   [1:0]                           m12_axi_gmem_RRESP,
    input                                   m12_axi_gmem_BVALID,
    output                                  m12_axi_gmem_BREADY,
    input   [1:0]                           m12_axi_gmem_BRESP,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m12_axi_gmem_BID,

    // AXI4 master interface 
    output                                  m13_axi_gmem_AWVALID,
    input                                   m13_axi_gmem_AWREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m13_axi_gmem_AWADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m13_axi_gmem_AWID,
    output  [7:0]                           m13_axi_gmem_AWLEN,
    output  [2:0]                           m13_axi_gmem_AWSIZE,
    output  [1:0]                           m13_axi_gmem_AWBURST,
    output  [1:0]                           m13_axi_gmem_AWLOCK,
    output  [3:0]                           m13_axi_gmem_AWCACHE,
    output  [2:0]                           m13_axi_gmem_AWPROT,
    output  [3:0]                           m13_axi_gmem_AWQOS,
    output  [3:0]                           m13_axi_gmem_AWREGION,
    output                                  m13_axi_gmem_WVALID,
    input                                   m13_axi_gmem_WREADY,
    output  [C_M_AXI_GMEM_DATA_WIDTH-1:0]   m13_axi_gmem_WDATA,
    output  [C_M_AXI_GMEM_DATA_WIDTH/8-1:0] m13_axi_gmem_WSTRB,
    output                                  m13_axi_gmem_WLAST,
    output                                  m13_axi_gmem_ARVALID,
    input                                   m13_axi_gmem_ARREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m13_axi_gmem_ARADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH-1:0]     m13_axi_gmem_ARID,
    output  [7:0]                           m13_axi_gmem_ARLEN,
    output  [2:0]                           m13_axi_gmem_ARSIZE,
    output  [1:0]                           m13_axi_gmem_ARBURST,
    output  [1:0]                           m13_axi_gmem_ARLOCK,
    output  [3:0]                           m13_axi_gmem_ARCACHE,
    output  [2:0]                           m13_axi_gmem_ARPROT,
    output  [3:0]                           m13_axi_gmem_ARQOS,
    output  [3:0]                           m13_axi_gmem_ARREGION,
    input                                   m13_axi_gmem_RVALID,
    output                                  m13_axi_gmem_RREADY,
    input   [C_M_AXI_GMEM_DATA_WIDTH - 1:0] m13_axi_gmem_RDATA,
    input                                   m13_axi_gmem_RLAST,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m13_axi_gmem_RID,
    input   [1:0]                           m13_axi_gmem_RRESP,
    input                                   m13_axi_gmem_BVALID,
    output                                  m13_axi_gmem_BREADY,
    input   [1:0]                           m13_axi_gmem_BRESP,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m13_axi_gmem_BID,

    // AXI4 master interface 
    output                                  m14_axi_gmem_AWVALID,
    input                                   m14_axi_gmem_AWREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m14_axi_gmem_AWADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m14_axi_gmem_AWID,
    output  [7:0]                           m14_axi_gmem_AWLEN,
    output  [2:0]                           m14_axi_gmem_AWSIZE,
    output  [1:0]                           m14_axi_gmem_AWBURST,
    output  [1:0]                           m14_axi_gmem_AWLOCK,
    output  [3:0]                           m14_axi_gmem_AWCACHE,
    output  [2:0]                           m14_axi_gmem_AWPROT,
    output  [3:0]                           m14_axi_gmem_AWQOS,
    output  [3:0]                           m14_axi_gmem_AWREGION,
    output                                  m14_axi_gmem_WVALID,
    input                                   m14_axi_gmem_WREADY,
    output  [C_M_AXI_GMEM_DATA_WIDTH-1:0]   m14_axi_gmem_WDATA,
    output  [C_M_AXI_GMEM_DATA_WIDTH/8-1:0] m14_axi_gmem_WSTRB,
    output                                  m14_axi_gmem_WLAST,
    output                                  m14_axi_gmem_ARVALID,
    input                                   m14_axi_gmem_ARREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m14_axi_gmem_ARADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH-1:0]     m14_axi_gmem_ARID,
    output  [7:0]                           m14_axi_gmem_ARLEN,
    output  [2:0]                           m14_axi_gmem_ARSIZE,
    output  [1:0]                           m14_axi_gmem_ARBURST,
    output  [1:0]                           m14_axi_gmem_ARLOCK,
    output  [3:0]                           m14_axi_gmem_ARCACHE,
    output  [2:0]                           m14_axi_gmem_ARPROT,
    output  [3:0]                           m14_axi_gmem_ARQOS,
    output  [3:0]                           m14_axi_gmem_ARREGION,
    input                                   m14_axi_gmem_RVALID,
    output                                  m14_axi_gmem_RREADY,
    input   [C_M_AXI_GMEM_DATA_WIDTH - 1:0] m14_axi_gmem_RDATA,
    input                                   m14_axi_gmem_RLAST,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m14_axi_gmem_RID,
    input   [1:0]                           m14_axi_gmem_RRESP,
    input                                   m14_axi_gmem_BVALID,
    output                                  m14_axi_gmem_BREADY,
    input   [1:0]                           m14_axi_gmem_BRESP,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m14_axi_gmem_BID,

    // AXI4 master interface 
    output                                  m15_axi_gmem_AWVALID,
    input                                   m15_axi_gmem_AWREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m15_axi_gmem_AWADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m15_axi_gmem_AWID,
    output  [7:0]                           m15_axi_gmem_AWLEN,
    output  [2:0]                           m15_axi_gmem_AWSIZE,
    output  [1:0]                           m15_axi_gmem_AWBURST,
    output  [1:0]                           m15_axi_gmem_AWLOCK,
    output  [3:0]                           m15_axi_gmem_AWCACHE,
    output  [2:0]                           m15_axi_gmem_AWPROT,
    output  [3:0]                           m15_axi_gmem_AWQOS,
    output  [3:0]                           m15_axi_gmem_AWREGION,
    output                                  m15_axi_gmem_WVALID,
    input                                   m15_axi_gmem_WREADY,
    output  [C_M_AXI_GMEM_DATA_WIDTH-1:0]   m15_axi_gmem_WDATA,
    output  [C_M_AXI_GMEM_DATA_WIDTH/8-1:0] m15_axi_gmem_WSTRB,
    output                                  m15_axi_gmem_WLAST,
    output                                  m15_axi_gmem_ARVALID,
    input                                   m15_axi_gmem_ARREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m15_axi_gmem_ARADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH-1:0]     m15_axi_gmem_ARID,
    output  [7:0]                           m15_axi_gmem_ARLEN,
    output  [2:0]                           m15_axi_gmem_ARSIZE,
    output  [1:0]                           m15_axi_gmem_ARBURST,
    output  [1:0]                           m15_axi_gmem_ARLOCK,
    output  [3:0]                           m15_axi_gmem_ARCACHE,
    output  [2:0]                           m15_axi_gmem_ARPROT,
    output  [3:0]                           m15_axi_gmem_ARQOS,
    output  [3:0]                           m15_axi_gmem_ARREGION,
    input                                   m15_axi_gmem_RVALID,
    output                                  m15_axi_gmem_RREADY,
    input   [C_M_AXI_GMEM_DATA_WIDTH - 1:0] m15_axi_gmem_RDATA,
    input                                   m15_axi_gmem_RLAST,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m15_axi_gmem_RID,
    input   [1:0]                           m15_axi_gmem_RRESP,
    input                                   m15_axi_gmem_BVALID,
    output                                  m15_axi_gmem_BREADY,
    input   [1:0]                           m15_axi_gmem_BRESP,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m15_axi_gmem_BID,

    // AXI4 master interface 
    output                                  m16_axi_gmem_AWVALID,
    input                                   m16_axi_gmem_AWREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m16_axi_gmem_AWADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m16_axi_gmem_AWID,
    output  [7:0]                           m16_axi_gmem_AWLEN,
    output  [2:0]                           m16_axi_gmem_AWSIZE,
    output  [1:0]                           m16_axi_gmem_AWBURST,
    output  [1:0]                           m16_axi_gmem_AWLOCK,
    output  [3:0]                           m16_axi_gmem_AWCACHE,
    output  [2:0]                           m16_axi_gmem_AWPROT,
    output  [3:0]                           m16_axi_gmem_AWQOS,
    output  [3:0]                           m16_axi_gmem_AWREGION,
    output                                  m16_axi_gmem_WVALID,
    input                                   m16_axi_gmem_WREADY,
    output  [C_M_AXI_GMEM_DATA_WIDTH-1:0]   m16_axi_gmem_WDATA,
    output  [C_M_AXI_GMEM_DATA_WIDTH/8-1:0] m16_axi_gmem_WSTRB,
    output                                  m16_axi_gmem_WLAST,
    output                                  m16_axi_gmem_ARVALID,
    input                                   m16_axi_gmem_ARREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m16_axi_gmem_ARADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH-1:0]     m16_axi_gmem_ARID,
    output  [7:0]                           m16_axi_gmem_ARLEN,
    output  [2:0]                           m16_axi_gmem_ARSIZE,
    output  [1:0]                           m16_axi_gmem_ARBURST,
    output  [1:0]                           m16_axi_gmem_ARLOCK,
    output  [3:0]                           m16_axi_gmem_ARCACHE,
    output  [2:0]                           m16_axi_gmem_ARPROT,
    output  [3:0]                           m16_axi_gmem_ARQOS,
    output  [3:0]                           m16_axi_gmem_ARREGION,
    input                                   m16_axi_gmem_RVALID,
    output                                  m16_axi_gmem_RREADY,
    input   [C_M_AXI_GMEM_DATA_WIDTH - 1:0] m16_axi_gmem_RDATA,
    input                                   m16_axi_gmem_RLAST,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m16_axi_gmem_RID,
    input   [1:0]                           m16_axi_gmem_RRESP,
    input                                   m16_axi_gmem_BVALID,
    output                                  m16_axi_gmem_BREADY,
    input   [1:0]                           m16_axi_gmem_BRESP,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m16_axi_gmem_BID,

    // AXI4 master interface 
    output                                  m17_axi_gmem_AWVALID,
    input                                   m17_axi_gmem_AWREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m17_axi_gmem_AWADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m17_axi_gmem_AWID,
    output  [7:0]                           m17_axi_gmem_AWLEN,
    output  [2:0]                           m17_axi_gmem_AWSIZE,
    output  [1:0]                           m17_axi_gmem_AWBURST,
    output  [1:0]                           m17_axi_gmem_AWLOCK,
    output  [3:0]                           m17_axi_gmem_AWCACHE,
    output  [2:0]                           m17_axi_gmem_AWPROT,
    output  [3:0]                           m17_axi_gmem_AWQOS,
    output  [3:0]                           m17_axi_gmem_AWREGION,
    output                                  m17_axi_gmem_WVALID,
    input                                   m17_axi_gmem_WREADY,
    output  [C_M_AXI_GMEM_DATA_WIDTH-1:0]   m17_axi_gmem_WDATA,
    output  [C_M_AXI_GMEM_DATA_WIDTH/8-1:0] m17_axi_gmem_WSTRB,
    output                                  m17_axi_gmem_WLAST,
    output                                  m17_axi_gmem_ARVALID,
    input                                   m17_axi_gmem_ARREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m17_axi_gmem_ARADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH-1:0]     m17_axi_gmem_ARID,
    output  [7:0]                           m17_axi_gmem_ARLEN,
    output  [2:0]                           m17_axi_gmem_ARSIZE,
    output  [1:0]                           m17_axi_gmem_ARBURST,
    output  [1:0]                           m17_axi_gmem_ARLOCK,
    output  [3:0]                           m17_axi_gmem_ARCACHE,
    output  [2:0]                           m17_axi_gmem_ARPROT,
    output  [3:0]                           m17_axi_gmem_ARQOS,
    output  [3:0]                           m17_axi_gmem_ARREGION,
    input                                   m17_axi_gmem_RVALID,
    output                                  m17_axi_gmem_RREADY,
    input   [C_M_AXI_GMEM_DATA_WIDTH - 1:0] m17_axi_gmem_RDATA,
    input                                   m17_axi_gmem_RLAST,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m17_axi_gmem_RID,
    input   [1:0]                           m17_axi_gmem_RRESP,
    input                                   m17_axi_gmem_BVALID,
    output                                  m17_axi_gmem_BREADY,
    input   [1:0]                           m17_axi_gmem_BRESP,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m17_axi_gmem_BID,

    // AXI4 master interface 
    output                                  m18_axi_gmem_AWVALID,
    input                                   m18_axi_gmem_AWREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m18_axi_gmem_AWADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m18_axi_gmem_AWID,
    output  [7:0]                           m18_axi_gmem_AWLEN,
    output  [2:0]                           m18_axi_gmem_AWSIZE,
    output  [1:0]                           m18_axi_gmem_AWBURST,
    output  [1:0]                           m18_axi_gmem_AWLOCK,
    output  [3:0]                           m18_axi_gmem_AWCACHE,
    output  [2:0]                           m18_axi_gmem_AWPROT,
    output  [3:0]                           m18_axi_gmem_AWQOS,
    output  [3:0]                           m18_axi_gmem_AWREGION,
    output                                  m18_axi_gmem_WVALID,
    input                                   m18_axi_gmem_WREADY,
    output  [C_M_AXI_GMEM_DATA_WIDTH-1:0]   m18_axi_gmem_WDATA,
    output  [C_M_AXI_GMEM_DATA_WIDTH/8-1:0] m18_axi_gmem_WSTRB,
    output                                  m18_axi_gmem_WLAST,
    output                                  m18_axi_gmem_ARVALID,
    input                                   m18_axi_gmem_ARREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m18_axi_gmem_ARADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH-1:0]     m18_axi_gmem_ARID,
    output  [7:0]                           m18_axi_gmem_ARLEN,
    output  [2:0]                           m18_axi_gmem_ARSIZE,
    output  [1:0]                           m18_axi_gmem_ARBURST,
    output  [1:0]                           m18_axi_gmem_ARLOCK,
    output  [3:0]                           m18_axi_gmem_ARCACHE,
    output  [2:0]                           m18_axi_gmem_ARPROT,
    output  [3:0]                           m18_axi_gmem_ARQOS,
    output  [3:0]                           m18_axi_gmem_ARREGION,
    input                                   m18_axi_gmem_RVALID,
    output                                  m18_axi_gmem_RREADY,
    input   [C_M_AXI_GMEM_DATA_WIDTH - 1:0] m18_axi_gmem_RDATA,
    input                                   m18_axi_gmem_RLAST,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m18_axi_gmem_RID,
    input   [1:0]                           m18_axi_gmem_RRESP,
    input                                   m18_axi_gmem_BVALID,
    output                                  m18_axi_gmem_BREADY,
    input   [1:0]                           m18_axi_gmem_BRESP,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m18_axi_gmem_BID,

    // AXI4 master interface 
    output                                  m19_axi_gmem_AWVALID,
    input                                   m19_axi_gmem_AWREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m19_axi_gmem_AWADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m19_axi_gmem_AWID,
    output  [7:0]                           m19_axi_gmem_AWLEN,
    output  [2:0]                           m19_axi_gmem_AWSIZE,
    output  [1:0]                           m19_axi_gmem_AWBURST,
    output  [1:0]                           m19_axi_gmem_AWLOCK,
    output  [3:0]                           m19_axi_gmem_AWCACHE,
    output  [2:0]                           m19_axi_gmem_AWPROT,
    output  [3:0]                           m19_axi_gmem_AWQOS,
    output  [3:0]                           m19_axi_gmem_AWREGION,
    output                                  m19_axi_gmem_WVALID,
    input                                   m19_axi_gmem_WREADY,
    output  [C_M_AXI_GMEM_DATA_WIDTH-1:0]   m19_axi_gmem_WDATA,
    output  [C_M_AXI_GMEM_DATA_WIDTH/8-1:0] m19_axi_gmem_WSTRB,
    output                                  m19_axi_gmem_WLAST,
    output                                  m19_axi_gmem_ARVALID,
    input                                   m19_axi_gmem_ARREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m19_axi_gmem_ARADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH-1:0]     m19_axi_gmem_ARID,
    output  [7:0]                           m19_axi_gmem_ARLEN,
    output  [2:0]                           m19_axi_gmem_ARSIZE,
    output  [1:0]                           m19_axi_gmem_ARBURST,
    output  [1:0]                           m19_axi_gmem_ARLOCK,
    output  [3:0]                           m19_axi_gmem_ARCACHE,
    output  [2:0]                           m19_axi_gmem_ARPROT,
    output  [3:0]                           m19_axi_gmem_ARQOS,
    output  [3:0]                           m19_axi_gmem_ARREGION,
    input                                   m19_axi_gmem_RVALID,
    output                                  m19_axi_gmem_RREADY,
    input   [C_M_AXI_GMEM_DATA_WIDTH - 1:0] m19_axi_gmem_RDATA,
    input                                   m19_axi_gmem_RLAST,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m19_axi_gmem_RID,
    input   [1:0]                           m19_axi_gmem_RRESP,
    input                                   m19_axi_gmem_BVALID,
    output                                  m19_axi_gmem_BREADY,
    input   [1:0]                           m19_axi_gmem_BRESP,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m19_axi_gmem_BID,

    // AXI4 master interface 
    output                                  m20_axi_gmem_AWVALID,
    input                                   m20_axi_gmem_AWREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m20_axi_gmem_AWADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m20_axi_gmem_AWID,
    output  [7:0]                           m20_axi_gmem_AWLEN,
    output  [2:0]                           m20_axi_gmem_AWSIZE,
    output  [1:0]                           m20_axi_gmem_AWBURST,
    output  [1:0]                           m20_axi_gmem_AWLOCK,
    output  [3:0]                           m20_axi_gmem_AWCACHE,
    output  [2:0]                           m20_axi_gmem_AWPROT,
    output  [3:0]                           m20_axi_gmem_AWQOS,
    output  [3:0]                           m20_axi_gmem_AWREGION,
    output                                  m20_axi_gmem_WVALID,
    input                                   m20_axi_gmem_WREADY,
    output  [C_M_AXI_GMEM_DATA_WIDTH-1:0]   m20_axi_gmem_WDATA,
    output  [C_M_AXI_GMEM_DATA_WIDTH/8-1:0] m20_axi_gmem_WSTRB,
    output                                  m20_axi_gmem_WLAST,
    output                                  m20_axi_gmem_ARVALID,
    input                                   m20_axi_gmem_ARREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m20_axi_gmem_ARADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH-1:0]     m20_axi_gmem_ARID,
    output  [7:0]                           m20_axi_gmem_ARLEN,
    output  [2:0]                           m20_axi_gmem_ARSIZE,
    output  [1:0]                           m20_axi_gmem_ARBURST,
    output  [1:0]                           m20_axi_gmem_ARLOCK,
    output  [3:0]                           m20_axi_gmem_ARCACHE,
    output  [2:0]                           m20_axi_gmem_ARPROT,
    output  [3:0]                           m20_axi_gmem_ARQOS,
    output  [3:0]                           m20_axi_gmem_ARREGION,
    input                                   m20_axi_gmem_RVALID,
    output                                  m20_axi_gmem_RREADY,
    input   [C_M_AXI_GMEM_DATA_WIDTH - 1:0] m20_axi_gmem_RDATA,
    input                                   m20_axi_gmem_RLAST,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m20_axi_gmem_RID,
    input   [1:0]                           m20_axi_gmem_RRESP,
    input                                   m20_axi_gmem_BVALID,
    output                                  m20_axi_gmem_BREADY,
    input   [1:0]                           m20_axi_gmem_BRESP,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m20_axi_gmem_BID,

    // AXI4 master interface 
    output                                  m21_axi_gmem_AWVALID,
    input                                   m21_axi_gmem_AWREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m21_axi_gmem_AWADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m21_axi_gmem_AWID,
    output  [7:0]                           m21_axi_gmem_AWLEN,
    output  [2:0]                           m21_axi_gmem_AWSIZE,
    output  [1:0]                           m21_axi_gmem_AWBURST,
    output  [1:0]                           m21_axi_gmem_AWLOCK,
    output  [3:0]                           m21_axi_gmem_AWCACHE,
    output  [2:0]                           m21_axi_gmem_AWPROT,
    output  [3:0]                           m21_axi_gmem_AWQOS,
    output  [3:0]                           m21_axi_gmem_AWREGION,
    output                                  m21_axi_gmem_WVALID,
    input                                   m21_axi_gmem_WREADY,
    output  [C_M_AXI_GMEM_DATA_WIDTH-1:0]   m21_axi_gmem_WDATA,
    output  [C_M_AXI_GMEM_DATA_WIDTH/8-1:0] m21_axi_gmem_WSTRB,
    output                                  m21_axi_gmem_WLAST,
    output                                  m21_axi_gmem_ARVALID,
    input                                   m21_axi_gmem_ARREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m21_axi_gmem_ARADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH-1:0]     m21_axi_gmem_ARID,
    output  [7:0]                           m21_axi_gmem_ARLEN,
    output  [2:0]                           m21_axi_gmem_ARSIZE,
    output  [1:0]                           m21_axi_gmem_ARBURST,
    output  [1:0]                           m21_axi_gmem_ARLOCK,
    output  [3:0]                           m21_axi_gmem_ARCACHE,
    output  [2:0]                           m21_axi_gmem_ARPROT,
    output  [3:0]                           m21_axi_gmem_ARQOS,
    output  [3:0]                           m21_axi_gmem_ARREGION,
    input                                   m21_axi_gmem_RVALID,
    output                                  m21_axi_gmem_RREADY,
    input   [C_M_AXI_GMEM_DATA_WIDTH - 1:0] m21_axi_gmem_RDATA,
    input                                   m21_axi_gmem_RLAST,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m21_axi_gmem_RID,
    input   [1:0]                           m21_axi_gmem_RRESP,
    input                                   m21_axi_gmem_BVALID,
    output                                  m21_axi_gmem_BREADY,
    input   [1:0]                           m21_axi_gmem_BRESP,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m21_axi_gmem_BID,

    // AXI4 master interface 
    output                                  m22_axi_gmem_AWVALID,
    input                                   m22_axi_gmem_AWREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m22_axi_gmem_AWADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m22_axi_gmem_AWID,
    output  [7:0]                           m22_axi_gmem_AWLEN,
    output  [2:0]                           m22_axi_gmem_AWSIZE,
    output  [1:0]                           m22_axi_gmem_AWBURST,
    output  [1:0]                           m22_axi_gmem_AWLOCK,
    output  [3:0]                           m22_axi_gmem_AWCACHE,
    output  [2:0]                           m22_axi_gmem_AWPROT,
    output  [3:0]                           m22_axi_gmem_AWQOS,
    output  [3:0]                           m22_axi_gmem_AWREGION,
    output                                  m22_axi_gmem_WVALID,
    input                                   m22_axi_gmem_WREADY,
    output  [C_M_AXI_GMEM_DATA_WIDTH-1:0]   m22_axi_gmem_WDATA,
    output  [C_M_AXI_GMEM_DATA_WIDTH/8-1:0] m22_axi_gmem_WSTRB,
    output                                  m22_axi_gmem_WLAST,
    output                                  m22_axi_gmem_ARVALID,
    input                                   m22_axi_gmem_ARREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m22_axi_gmem_ARADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH-1:0]     m22_axi_gmem_ARID,
    output  [7:0]                           m22_axi_gmem_ARLEN,
    output  [2:0]                           m22_axi_gmem_ARSIZE,
    output  [1:0]                           m22_axi_gmem_ARBURST,
    output  [1:0]                           m22_axi_gmem_ARLOCK,
    output  [3:0]                           m22_axi_gmem_ARCACHE,
    output  [2:0]                           m22_axi_gmem_ARPROT,
    output  [3:0]                           m22_axi_gmem_ARQOS,
    output  [3:0]                           m22_axi_gmem_ARREGION,
    input                                   m22_axi_gmem_RVALID,
    output                                  m22_axi_gmem_RREADY,
    input   [C_M_AXI_GMEM_DATA_WIDTH - 1:0] m22_axi_gmem_RDATA,
    input                                   m22_axi_gmem_RLAST,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m22_axi_gmem_RID,
    input   [1:0]                           m22_axi_gmem_RRESP,
    input                                   m22_axi_gmem_BVALID,
    output                                  m22_axi_gmem_BREADY,
    input   [1:0]                           m22_axi_gmem_BRESP,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m22_axi_gmem_BID,

    // AXI4 master interface 
    output                                  m23_axi_gmem_AWVALID,
    input                                   m23_axi_gmem_AWREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m23_axi_gmem_AWADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m23_axi_gmem_AWID,
    output  [7:0]                           m23_axi_gmem_AWLEN,
    output  [2:0]                           m23_axi_gmem_AWSIZE,
    output  [1:0]                           m23_axi_gmem_AWBURST,
    output  [1:0]                           m23_axi_gmem_AWLOCK,
    output  [3:0]                           m23_axi_gmem_AWCACHE,
    output  [2:0]                           m23_axi_gmem_AWPROT,
    output  [3:0]                           m23_axi_gmem_AWQOS,
    output  [3:0]                           m23_axi_gmem_AWREGION,
    output                                  m23_axi_gmem_WVALID,
    input                                   m23_axi_gmem_WREADY,
    output  [C_M_AXI_GMEM_DATA_WIDTH-1:0]   m23_axi_gmem_WDATA,
    output  [C_M_AXI_GMEM_DATA_WIDTH/8-1:0] m23_axi_gmem_WSTRB,
    output                                  m23_axi_gmem_WLAST,
    output                                  m23_axi_gmem_ARVALID,
    input                                   m23_axi_gmem_ARREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m23_axi_gmem_ARADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH-1:0]     m23_axi_gmem_ARID,
    output  [7:0]                           m23_axi_gmem_ARLEN,
    output  [2:0]                           m23_axi_gmem_ARSIZE,
    output  [1:0]                           m23_axi_gmem_ARBURST,
    output  [1:0]                           m23_axi_gmem_ARLOCK,
    output  [3:0]                           m23_axi_gmem_ARCACHE,
    output  [2:0]                           m23_axi_gmem_ARPROT,
    output  [3:0]                           m23_axi_gmem_ARQOS,
    output  [3:0]                           m23_axi_gmem_ARREGION,
    input                                   m23_axi_gmem_RVALID,
    output                                  m23_axi_gmem_RREADY,
    input   [C_M_AXI_GMEM_DATA_WIDTH - 1:0] m23_axi_gmem_RDATA,
    input                                   m23_axi_gmem_RLAST,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m23_axi_gmem_RID,
    input   [1:0]                           m23_axi_gmem_RRESP,
    input                                   m23_axi_gmem_BVALID,
    output                                  m23_axi_gmem_BREADY,
    input   [1:0]                           m23_axi_gmem_BRESP,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m23_axi_gmem_BID,

    // AXI4 master interface 
    output                                  m24_axi_gmem_AWVALID,
    input                                   m24_axi_gmem_AWREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m24_axi_gmem_AWADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m24_axi_gmem_AWID,
    output  [7:0]                           m24_axi_gmem_AWLEN,
    output  [2:0]                           m24_axi_gmem_AWSIZE,
    output  [1:0]                           m24_axi_gmem_AWBURST,
    output  [1:0]                           m24_axi_gmem_AWLOCK,
    output  [3:0]                           m24_axi_gmem_AWCACHE,
    output  [2:0]                           m24_axi_gmem_AWPROT,
    output  [3:0]                           m24_axi_gmem_AWQOS,
    output  [3:0]                           m24_axi_gmem_AWREGION,
    output                                  m24_axi_gmem_WVALID,
    input                                   m24_axi_gmem_WREADY,
    output  [C_M_AXI_GMEM_DATA_WIDTH-1:0]   m24_axi_gmem_WDATA,
    output  [C_M_AXI_GMEM_DATA_WIDTH/8-1:0] m24_axi_gmem_WSTRB,
    output                                  m24_axi_gmem_WLAST,
    output                                  m24_axi_gmem_ARVALID,
    input                                   m24_axi_gmem_ARREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m24_axi_gmem_ARADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH-1:0]     m24_axi_gmem_ARID,
    output  [7:0]                           m24_axi_gmem_ARLEN,
    output  [2:0]                           m24_axi_gmem_ARSIZE,
    output  [1:0]                           m24_axi_gmem_ARBURST,
    output  [1:0]                           m24_axi_gmem_ARLOCK,
    output  [3:0]                           m24_axi_gmem_ARCACHE,
    output  [2:0]                           m24_axi_gmem_ARPROT,
    output  [3:0]                           m24_axi_gmem_ARQOS,
    output  [3:0]                           m24_axi_gmem_ARREGION,
    input                                   m24_axi_gmem_RVALID,
    output                                  m24_axi_gmem_RREADY,
    input   [C_M_AXI_GMEM_DATA_WIDTH - 1:0] m24_axi_gmem_RDATA,
    input                                   m24_axi_gmem_RLAST,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m24_axi_gmem_RID,
    input   [1:0]                           m24_axi_gmem_RRESP,
    input                                   m24_axi_gmem_BVALID,
    output                                  m24_axi_gmem_BREADY,
    input   [1:0]                           m24_axi_gmem_BRESP,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m24_axi_gmem_BID,

    // AXI4 master interface 
    output                                  m25_axi_gmem_AWVALID,
    input                                   m25_axi_gmem_AWREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m25_axi_gmem_AWADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m25_axi_gmem_AWID,
    output  [7:0]                           m25_axi_gmem_AWLEN,
    output  [2:0]                           m25_axi_gmem_AWSIZE,
    output  [1:0]                           m25_axi_gmem_AWBURST,
    output  [1:0]                           m25_axi_gmem_AWLOCK,
    output  [3:0]                           m25_axi_gmem_AWCACHE,
    output  [2:0]                           m25_axi_gmem_AWPROT,
    output  [3:0]                           m25_axi_gmem_AWQOS,
    output  [3:0]                           m25_axi_gmem_AWREGION,
    output                                  m25_axi_gmem_WVALID,
    input                                   m25_axi_gmem_WREADY,
    output  [C_M_AXI_GMEM_DATA_WIDTH-1:0]   m25_axi_gmem_WDATA,
    output  [C_M_AXI_GMEM_DATA_WIDTH/8-1:0] m25_axi_gmem_WSTRB,
    output                                  m25_axi_gmem_WLAST,
    output                                  m25_axi_gmem_ARVALID,
    input                                   m25_axi_gmem_ARREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m25_axi_gmem_ARADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH-1:0]     m25_axi_gmem_ARID,
    output  [7:0]                           m25_axi_gmem_ARLEN,
    output  [2:0]                           m25_axi_gmem_ARSIZE,
    output  [1:0]                           m25_axi_gmem_ARBURST,
    output  [1:0]                           m25_axi_gmem_ARLOCK,
    output  [3:0]                           m25_axi_gmem_ARCACHE,
    output  [2:0]                           m25_axi_gmem_ARPROT,
    output  [3:0]                           m25_axi_gmem_ARQOS,
    output  [3:0]                           m25_axi_gmem_ARREGION,
    input                                   m25_axi_gmem_RVALID,
    output                                  m25_axi_gmem_RREADY,
    input   [C_M_AXI_GMEM_DATA_WIDTH - 1:0] m25_axi_gmem_RDATA,
    input                                   m25_axi_gmem_RLAST,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m25_axi_gmem_RID,
    input   [1:0]                           m25_axi_gmem_RRESP,
    input                                   m25_axi_gmem_BVALID,
    output                                  m25_axi_gmem_BREADY,
    input   [1:0]                           m25_axi_gmem_BRESP,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m25_axi_gmem_BID,

    // AXI4 master interface 
    output                                  m26_axi_gmem_AWVALID,
    input                                   m26_axi_gmem_AWREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m26_axi_gmem_AWADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m26_axi_gmem_AWID,
    output  [7:0]                           m26_axi_gmem_AWLEN,
    output  [2:0]                           m26_axi_gmem_AWSIZE,
    output  [1:0]                           m26_axi_gmem_AWBURST,
    output  [1:0]                           m26_axi_gmem_AWLOCK,
    output  [3:0]                           m26_axi_gmem_AWCACHE,
    output  [2:0]                           m26_axi_gmem_AWPROT,
    output  [3:0]                           m26_axi_gmem_AWQOS,
    output  [3:0]                           m26_axi_gmem_AWREGION,
    output                                  m26_axi_gmem_WVALID,
    input                                   m26_axi_gmem_WREADY,
    output  [C_M_AXI_GMEM_DATA_WIDTH-1:0]   m26_axi_gmem_WDATA,
    output  [C_M_AXI_GMEM_DATA_WIDTH/8-1:0] m26_axi_gmem_WSTRB,
    output                                  m26_axi_gmem_WLAST,
    output                                  m26_axi_gmem_ARVALID,
    input                                   m26_axi_gmem_ARREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m26_axi_gmem_ARADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH-1:0]     m26_axi_gmem_ARID,
    output  [7:0]                           m26_axi_gmem_ARLEN,
    output  [2:0]                           m26_axi_gmem_ARSIZE,
    output  [1:0]                           m26_axi_gmem_ARBURST,
    output  [1:0]                           m26_axi_gmem_ARLOCK,
    output  [3:0]                           m26_axi_gmem_ARCACHE,
    output  [2:0]                           m26_axi_gmem_ARPROT,
    output  [3:0]                           m26_axi_gmem_ARQOS,
    output  [3:0]                           m26_axi_gmem_ARREGION,
    input                                   m26_axi_gmem_RVALID,
    output                                  m26_axi_gmem_RREADY,
    input   [C_M_AXI_GMEM_DATA_WIDTH - 1:0] m26_axi_gmem_RDATA,
    input                                   m26_axi_gmem_RLAST,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m26_axi_gmem_RID,
    input   [1:0]                           m26_axi_gmem_RRESP,
    input                                   m26_axi_gmem_BVALID,
    output                                  m26_axi_gmem_BREADY,
    input   [1:0]                           m26_axi_gmem_BRESP,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m26_axi_gmem_BID,

    // AXI4 master interface 
    output                                  m27_axi_gmem_AWVALID,
    input                                   m27_axi_gmem_AWREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m27_axi_gmem_AWADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m27_axi_gmem_AWID,
    output  [7:0]                           m27_axi_gmem_AWLEN,
    output  [2:0]                           m27_axi_gmem_AWSIZE,
    output  [1:0]                           m27_axi_gmem_AWBURST,
    output  [1:0]                           m27_axi_gmem_AWLOCK,
    output  [3:0]                           m27_axi_gmem_AWCACHE,
    output  [2:0]                           m27_axi_gmem_AWPROT,
    output  [3:0]                           m27_axi_gmem_AWQOS,
    output  [3:0]                           m27_axi_gmem_AWREGION,
    output                                  m27_axi_gmem_WVALID,
    input                                   m27_axi_gmem_WREADY,
    output  [C_M_AXI_GMEM_DATA_WIDTH-1:0]   m27_axi_gmem_WDATA,
    output  [C_M_AXI_GMEM_DATA_WIDTH/8-1:0] m27_axi_gmem_WSTRB,
    output                                  m27_axi_gmem_WLAST,
    output                                  m27_axi_gmem_ARVALID,
    input                                   m27_axi_gmem_ARREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m27_axi_gmem_ARADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH-1:0]     m27_axi_gmem_ARID,
    output  [7:0]                           m27_axi_gmem_ARLEN,
    output  [2:0]                           m27_axi_gmem_ARSIZE,
    output  [1:0]                           m27_axi_gmem_ARBURST,
    output  [1:0]                           m27_axi_gmem_ARLOCK,
    output  [3:0]                           m27_axi_gmem_ARCACHE,
    output  [2:0]                           m27_axi_gmem_ARPROT,
    output  [3:0]                           m27_axi_gmem_ARQOS,
    output  [3:0]                           m27_axi_gmem_ARREGION,
    input                                   m27_axi_gmem_RVALID,
    output                                  m27_axi_gmem_RREADY,
    input   [C_M_AXI_GMEM_DATA_WIDTH - 1:0] m27_axi_gmem_RDATA,
    input                                   m27_axi_gmem_RLAST,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m27_axi_gmem_RID,
    input   [1:0]                           m27_axi_gmem_RRESP,
    input                                   m27_axi_gmem_BVALID,
    output                                  m27_axi_gmem_BREADY,
    input   [1:0]                           m27_axi_gmem_BRESP,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m27_axi_gmem_BID,

    // AXI4 master interface 
    output                                  m28_axi_gmem_AWVALID,
    input                                   m28_axi_gmem_AWREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m28_axi_gmem_AWADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m28_axi_gmem_AWID,
    output  [7:0]                           m28_axi_gmem_AWLEN,
    output  [2:0]                           m28_axi_gmem_AWSIZE,
    output  [1:0]                           m28_axi_gmem_AWBURST,
    output  [1:0]                           m28_axi_gmem_AWLOCK,
    output  [3:0]                           m28_axi_gmem_AWCACHE,
    output  [2:0]                           m28_axi_gmem_AWPROT,
    output  [3:0]                           m28_axi_gmem_AWQOS,
    output  [3:0]                           m28_axi_gmem_AWREGION,
    output                                  m28_axi_gmem_WVALID,
    input                                   m28_axi_gmem_WREADY,
    output  [C_M_AXI_GMEM_DATA_WIDTH-1:0]   m28_axi_gmem_WDATA,
    output  [C_M_AXI_GMEM_DATA_WIDTH/8-1:0] m28_axi_gmem_WSTRB,
    output                                  m28_axi_gmem_WLAST,
    output                                  m28_axi_gmem_ARVALID,
    input                                   m28_axi_gmem_ARREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m28_axi_gmem_ARADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH-1:0]     m28_axi_gmem_ARID,
    output  [7:0]                           m28_axi_gmem_ARLEN,
    output  [2:0]                           m28_axi_gmem_ARSIZE,
    output  [1:0]                           m28_axi_gmem_ARBURST,
    output  [1:0]                           m28_axi_gmem_ARLOCK,
    output  [3:0]                           m28_axi_gmem_ARCACHE,
    output  [2:0]                           m28_axi_gmem_ARPROT,
    output  [3:0]                           m28_axi_gmem_ARQOS,
    output  [3:0]                           m28_axi_gmem_ARREGION,
    input                                   m28_axi_gmem_RVALID,
    output                                  m28_axi_gmem_RREADY,
    input   [C_M_AXI_GMEM_DATA_WIDTH - 1:0] m28_axi_gmem_RDATA,
    input                                   m28_axi_gmem_RLAST,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m28_axi_gmem_RID,
    input   [1:0]                           m28_axi_gmem_RRESP,
    input                                   m28_axi_gmem_BVALID,
    output                                  m28_axi_gmem_BREADY,
    input   [1:0]                           m28_axi_gmem_BRESP,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m28_axi_gmem_BID,

    // AXI4 master interface 
    output                                  m29_axi_gmem_AWVALID,
    input                                   m29_axi_gmem_AWREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m29_axi_gmem_AWADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m29_axi_gmem_AWID,
    output  [7:0]                           m29_axi_gmem_AWLEN,
    output  [2:0]                           m29_axi_gmem_AWSIZE,
    output  [1:0]                           m29_axi_gmem_AWBURST,
    output  [1:0]                           m29_axi_gmem_AWLOCK,
    output  [3:0]                           m29_axi_gmem_AWCACHE,
    output  [2:0]                           m29_axi_gmem_AWPROT,
    output  [3:0]                           m29_axi_gmem_AWQOS,
    output  [3:0]                           m29_axi_gmem_AWREGION,
    output                                  m29_axi_gmem_WVALID,
    input                                   m29_axi_gmem_WREADY,
    output  [C_M_AXI_GMEM_DATA_WIDTH-1:0]   m29_axi_gmem_WDATA,
    output  [C_M_AXI_GMEM_DATA_WIDTH/8-1:0] m29_axi_gmem_WSTRB,
    output                                  m29_axi_gmem_WLAST,
    output                                  m29_axi_gmem_ARVALID,
    input                                   m29_axi_gmem_ARREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m29_axi_gmem_ARADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH-1:0]     m29_axi_gmem_ARID,
    output  [7:0]                           m29_axi_gmem_ARLEN,
    output  [2:0]                           m29_axi_gmem_ARSIZE,
    output  [1:0]                           m29_axi_gmem_ARBURST,
    output  [1:0]                           m29_axi_gmem_ARLOCK,
    output  [3:0]                           m29_axi_gmem_ARCACHE,
    output  [2:0]                           m29_axi_gmem_ARPROT,
    output  [3:0]                           m29_axi_gmem_ARQOS,
    output  [3:0]                           m29_axi_gmem_ARREGION,
    input                                   m29_axi_gmem_RVALID,
    output                                  m29_axi_gmem_RREADY,
    input   [C_M_AXI_GMEM_DATA_WIDTH - 1:0] m29_axi_gmem_RDATA,
    input                                   m29_axi_gmem_RLAST,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m29_axi_gmem_RID,
    input   [1:0]                           m29_axi_gmem_RRESP,
    input                                   m29_axi_gmem_BVALID,
    output                                  m29_axi_gmem_BREADY,
    input   [1:0]                           m29_axi_gmem_BRESP,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m29_axi_gmem_BID,

    // AXI4 master interface 
    output                                  m30_axi_gmem_AWVALID,
    input                                   m30_axi_gmem_AWREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m30_axi_gmem_AWADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m30_axi_gmem_AWID,
    output  [7:0]                           m30_axi_gmem_AWLEN,
    output  [2:0]                           m30_axi_gmem_AWSIZE,
    output  [1:0]                           m30_axi_gmem_AWBURST,
    output  [1:0]                           m30_axi_gmem_AWLOCK,
    output  [3:0]                           m30_axi_gmem_AWCACHE,
    output  [2:0]                           m30_axi_gmem_AWPROT,
    output  [3:0]                           m30_axi_gmem_AWQOS,
    output  [3:0]                           m30_axi_gmem_AWREGION,
    output                                  m30_axi_gmem_WVALID,
    input                                   m30_axi_gmem_WREADY,
    output  [C_M_AXI_GMEM_DATA_WIDTH-1:0]   m30_axi_gmem_WDATA,
    output  [C_M_AXI_GMEM_DATA_WIDTH/8-1:0] m30_axi_gmem_WSTRB,
    output                                  m30_axi_gmem_WLAST,
    output                                  m30_axi_gmem_ARVALID,
    input                                   m30_axi_gmem_ARREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m30_axi_gmem_ARADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH-1:0]     m30_axi_gmem_ARID,
    output  [7:0]                           m30_axi_gmem_ARLEN,
    output  [2:0]                           m30_axi_gmem_ARSIZE,
    output  [1:0]                           m30_axi_gmem_ARBURST,
    output  [1:0]                           m30_axi_gmem_ARLOCK,
    output  [3:0]                           m30_axi_gmem_ARCACHE,
    output  [2:0]                           m30_axi_gmem_ARPROT,
    output  [3:0]                           m30_axi_gmem_ARQOS,
    output  [3:0]                           m30_axi_gmem_ARREGION,
    input                                   m30_axi_gmem_RVALID,
    output                                  m30_axi_gmem_RREADY,
    input   [C_M_AXI_GMEM_DATA_WIDTH - 1:0] m30_axi_gmem_RDATA,
    input                                   m30_axi_gmem_RLAST,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m30_axi_gmem_RID,
    input   [1:0]                           m30_axi_gmem_RRESP,
    input                                   m30_axi_gmem_BVALID,
    output                                  m30_axi_gmem_BREADY,
    input   [1:0]                           m30_axi_gmem_BRESP,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m30_axi_gmem_BID,

    // AXI4 master interface 
    output                                  m31_axi_gmem_AWVALID,
    input                                   m31_axi_gmem_AWREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m31_axi_gmem_AWADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m31_axi_gmem_AWID,
    output  [7:0]                           m31_axi_gmem_AWLEN,
    output  [2:0]                           m31_axi_gmem_AWSIZE,
    output  [1:0]                           m31_axi_gmem_AWBURST,
    output  [1:0]                           m31_axi_gmem_AWLOCK,
    output  [3:0]                           m31_axi_gmem_AWCACHE,
    output  [2:0]                           m31_axi_gmem_AWPROT,
    output  [3:0]                           m31_axi_gmem_AWQOS,
    output  [3:0]                           m31_axi_gmem_AWREGION,
    output                                  m31_axi_gmem_WVALID,
    input                                   m31_axi_gmem_WREADY,
    output  [C_M_AXI_GMEM_DATA_WIDTH-1:0]   m31_axi_gmem_WDATA,
    output  [C_M_AXI_GMEM_DATA_WIDTH/8-1:0] m31_axi_gmem_WSTRB,
    output                                  m31_axi_gmem_WLAST,
    output                                  m31_axi_gmem_ARVALID,
    input                                   m31_axi_gmem_ARREADY,
    output  [C_M_AXI_GMEM_ADDR_WIDTH-1:0]   m31_axi_gmem_ARADDR,
    output  [C_M_AXI_GMEM_ID_WIDTH-1:0]     m31_axi_gmem_ARID,
    output  [7:0]                           m31_axi_gmem_ARLEN,
    output  [2:0]                           m31_axi_gmem_ARSIZE,
    output  [1:0]                           m31_axi_gmem_ARBURST,
    output  [1:0]                           m31_axi_gmem_ARLOCK,
    output  [3:0]                           m31_axi_gmem_ARCACHE,
    output  [2:0]                           m31_axi_gmem_ARPROT,
    output  [3:0]                           m31_axi_gmem_ARQOS,
    output  [3:0]                           m31_axi_gmem_ARREGION,
    input                                   m31_axi_gmem_RVALID,
    output                                  m31_axi_gmem_RREADY,
    input   [C_M_AXI_GMEM_DATA_WIDTH - 1:0] m31_axi_gmem_RDATA,
    input                                   m31_axi_gmem_RLAST,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m31_axi_gmem_RID,
    input   [1:0]                           m31_axi_gmem_RRESP,
    input                                   m31_axi_gmem_BVALID,
    output                                  m31_axi_gmem_BREADY,
    input   [1:0]                           m31_axi_gmem_BRESP,
    input   [C_M_AXI_GMEM_ID_WIDTH - 1:0]   m31_axi_gmem_BID,

    // AXI4-Lite slave interface
    input  wire                                    s_axi_control_AWVALID,
    output wire                                    s_axi_control_AWREADY,
    input  wire [C_S_AXI_CONTROL_ADDR_WIDTH-1:0]   s_axi_control_AWADDR,
    input  wire                                    s_axi_control_WVALID,
    output wire                                    s_axi_control_WREADY,
    input  wire [C_S_AXI_CONTROL_DATA_WIDTH-1:0]   s_axi_control_WDATA,
    input  wire [C_S_AXI_CONTROL_DATA_WIDTH/8-1:0] s_axi_control_WSTRB,
    input  wire                                    s_axi_control_ARVALID,
    output wire                                    s_axi_control_ARREADY,
    input  wire [C_S_AXI_CONTROL_ADDR_WIDTH-1:0]   s_axi_control_ARADDR,
    output wire                                    s_axi_control_RVALID,
    input  wire                                    s_axi_control_RREADY,
    output wire [C_S_AXI_CONTROL_DATA_WIDTH-1:0]   s_axi_control_RDATA,
    output wire [1:0]                              s_axi_control_RRESP,
    output wire                                    s_axi_control_BVALID,
    input  wire                                    s_axi_control_BREADY,
    output wire [1:0]                              s_axi_control_BRESP,
    output wire                                    interrupt
);
    ///////////////////////////////////////////////////////////////////////////////
    // Local Parameters (constants)
    ///////////////////////////////////////////////////////////////////////////////
    localparam integer LP_NUM_READ_CHANNELS  = 2;
    localparam integer LP_LENGTH_WIDTH       = 32;
    localparam integer LP_DW_BYTES           = C_M_AXI_GMEM_DATA_WIDTH/8;
    localparam integer LP_AXI_BURST_LEN      = 4096/LP_DW_BYTES < 256 ? 4096/LP_DW_BYTES : 256;
    localparam integer LP_LOG_BURST_LEN      = $clog2(LP_AXI_BURST_LEN);
    localparam integer LP_RD_MAX_OUTSTANDING = 3;
    localparam integer LP_RD_FIFO_DEPTH      = LP_AXI_BURST_LEN*(LP_RD_MAX_OUTSTANDING + 1);
    localparam integer LP_WR_FIFO_DEPTH      = LP_AXI_BURST_LEN;

    ///////////////////////////////////////////////////////////////////////////////
    // Variables
    ///////////////////////////////////////////////////////////////////////////////
    wire ap_start;
    wire ap_start_pulse;
    wire ap_ready;
    wire ap_done;
    reg areset = 1'b0;
    reg ap_idle = 1'b1;
    reg ap_start_r;

    wire dev_reset;
    wire dev_continue;
    wire [1:0] dev_bytemode;
    wire dev_done;
    wire dev_start;
    wire dev_load_text;
    
    wire key_first;
    wire key_begingap;
    wire key_endgap;
    wire key_last;
    wire key_mask;
    wire [1:0]key_bytemode;
    wire [7:0]key_data;
    wire [5:0]key_len;

    wire result_rden;
    wire [15:0] result_data;
    wire result_valid;
    wire [31:0] bash_code;

    wire bitstream_rden;
    wire [63:0]bitstream;
    wire [31:0]match_count;
    wire match_count_vld;

    wire [31:0]ikey;
    wire ikey_wren;

    wire [31:0]                rd_done;
    wire [31:0]                rd_done2;
    wire [63:0]                rd_addr  [0:31];
    wire [31:0]                rd_length[0:31];
    wire [31:0]                rd_en;
    wire [63:0]                rd_data  [0:31];
    wire [31:0]                rd_datavld;
    wire [31:0]                rd_tvalid_n;

    wire [63:0] start_addr;
    wire [63:0] file_size;
    wire [31:0] load_start;

    wire                       ctrl_load_filesize;
    wire                       ctrl_load_address;
    wire [63:0]                fm_next_filesize;
    wire [63:0]                fm_next_address;
    wire                       fm_overlap;
    wire                       fm_done;
    wire                       fm_ready;
    wire [63:0]                fm_bash_offset;
    wire [31:0]                fm_bashcount;
    wire                       fm_bashupdate;
    
    wire [31:0] count0;
    wire [31:0] count1;
    wire [31:0] rd_channel_idle;
    ///////////////////////////////////////////////////////////////////////////////
    // RTL Logic 
    ///////////////////////////////////////////////////////////////////////////////
    // Tie-off unused AXI protocol features
    assign m00_axi_gmem_AWID     = {C_M_AXI_GMEM_ID_WIDTH{1'b0}};
    assign m00_axi_gmem_AWBURST  = 2'b01;
    assign m00_axi_gmem_AWLOCK   = 2'b00;
    assign m00_axi_gmem_AWCACHE  = 4'b0011;
    assign m00_axi_gmem_AWPROT   = 3'b000;
    assign m00_axi_gmem_AWQOS    = 4'b0000;
    assign m00_axi_gmem_AWREGION = 4'b0000;
    assign m00_axi_gmem_ARBURST  = 2'b01;
    assign m00_axi_gmem_ARLOCK   = 2'b00;
    assign m00_axi_gmem_ARCACHE  = 4'b0011;
    assign m00_axi_gmem_ARPROT   = 3'b000;
    assign m00_axi_gmem_ARQOS    = 4'b0000;
    assign m00_axi_gmem_ARREGION = 4'b0000;

    assign m01_axi_gmem_AWID     = {C_M_AXI_GMEM_ID_WIDTH{1'b0}};
    assign m01_axi_gmem_AWBURST  = 2'b01;
    assign m01_axi_gmem_AWLOCK   = 2'b00;
    assign m01_axi_gmem_AWCACHE  = 4'b0011;
    assign m01_axi_gmem_AWPROT   = 3'b000;
    assign m01_axi_gmem_AWQOS    = 4'b0000;
    assign m01_axi_gmem_AWREGION = 4'b0000;
    assign m01_axi_gmem_ARBURST  = 2'b01;
    assign m01_axi_gmem_ARLOCK   = 2'b00;
    assign m01_axi_gmem_ARCACHE  = 4'b0011;
    assign m01_axi_gmem_ARPROT   = 3'b000;
    assign m01_axi_gmem_ARQOS    = 4'b0000;
    assign m01_axi_gmem_ARREGION = 4'b0000;

    assign m02_axi_gmem_AWID     = {C_M_AXI_GMEM_ID_WIDTH{1'b0}};
    assign m02_axi_gmem_AWBURST  = 2'b01;
    assign m02_axi_gmem_AWLOCK   = 2'b00;
    assign m02_axi_gmem_AWCACHE  = 4'b0011;
    assign m02_axi_gmem_AWPROT   = 3'b000;
    assign m02_axi_gmem_AWQOS    = 4'b0000;
    assign m02_axi_gmem_AWREGION = 4'b0000;
    assign m02_axi_gmem_ARBURST  = 2'b01;
    assign m02_axi_gmem_ARLOCK   = 2'b00;
    assign m02_axi_gmem_ARCACHE  = 4'b0011;
    assign m02_axi_gmem_ARPROT   = 3'b000;
    assign m02_axi_gmem_ARQOS    = 4'b0000;
    assign m02_axi_gmem_ARREGION = 4'b0000;

    assign m03_axi_gmem_AWID     = {C_M_AXI_GMEM_ID_WIDTH{1'b0}};
    assign m03_axi_gmem_AWBURST  = 2'b01;
    assign m03_axi_gmem_AWLOCK   = 2'b00;
    assign m03_axi_gmem_AWCACHE  = 4'b0011;
    assign m03_axi_gmem_AWPROT   = 3'b000;
    assign m03_axi_gmem_AWQOS    = 4'b0000;
    assign m03_axi_gmem_AWREGION = 4'b0000;
    assign m03_axi_gmem_ARBURST  = 2'b01;
    assign m03_axi_gmem_ARLOCK   = 2'b00;
    assign m03_axi_gmem_ARCACHE  = 4'b0011;
    assign m03_axi_gmem_ARPROT   = 3'b000;
    assign m03_axi_gmem_ARQOS    = 4'b0000;
    assign m03_axi_gmem_ARREGION = 4'b0000;

    assign m04_axi_gmem_AWID     = {C_M_AXI_GMEM_ID_WIDTH{1'b0}};
    assign m04_axi_gmem_AWBURST  = 2'b01;
    assign m04_axi_gmem_AWLOCK   = 2'b00;
    assign m04_axi_gmem_AWCACHE  = 4'b0011;
    assign m04_axi_gmem_AWPROT   = 3'b000;
    assign m04_axi_gmem_AWQOS    = 4'b0000;
    assign m04_axi_gmem_AWREGION = 4'b0000;
    assign m04_axi_gmem_ARBURST  = 2'b01;
    assign m04_axi_gmem_ARLOCK   = 2'b00;
    assign m04_axi_gmem_ARCACHE  = 4'b0011;
    assign m04_axi_gmem_ARPROT   = 3'b000;
    assign m04_axi_gmem_ARQOS    = 4'b0000;
    assign m04_axi_gmem_ARREGION = 4'b0000;

    assign m05_axi_gmem_AWID     = {C_M_AXI_GMEM_ID_WIDTH{1'b0}};
    assign m05_axi_gmem_AWBURST  = 2'b01;
    assign m05_axi_gmem_AWLOCK   = 2'b00;
    assign m05_axi_gmem_AWCACHE  = 4'b0011;
    assign m05_axi_gmem_AWPROT   = 3'b000;
    assign m05_axi_gmem_AWQOS    = 4'b0000;
    assign m05_axi_gmem_AWREGION = 4'b0000;
    assign m05_axi_gmem_ARBURST  = 2'b01;
    assign m05_axi_gmem_ARLOCK   = 2'b00;
    assign m05_axi_gmem_ARCACHE  = 4'b0011;
    assign m05_axi_gmem_ARPROT   = 3'b000;
    assign m05_axi_gmem_ARQOS    = 4'b0000;
    assign m05_axi_gmem_ARREGION = 4'b0000;

    assign m06_axi_gmem_AWID     = {C_M_AXI_GMEM_ID_WIDTH{1'b0}};
    assign m06_axi_gmem_AWBURST  = 2'b01;
    assign m06_axi_gmem_AWLOCK   = 2'b00;
    assign m06_axi_gmem_AWCACHE  = 4'b0011;
    assign m06_axi_gmem_AWPROT   = 3'b000;
    assign m06_axi_gmem_AWQOS    = 4'b0000;
    assign m06_axi_gmem_AWREGION = 4'b0000;
    assign m06_axi_gmem_ARBURST  = 2'b01;
    assign m06_axi_gmem_ARLOCK   = 2'b00;
    assign m06_axi_gmem_ARCACHE  = 4'b0011;
    assign m06_axi_gmem_ARPROT   = 3'b000;
    assign m06_axi_gmem_ARQOS    = 4'b0000;
    assign m06_axi_gmem_ARREGION = 4'b0000;

    assign m07_axi_gmem_AWID     = {C_M_AXI_GMEM_ID_WIDTH{1'b0}};
    assign m07_axi_gmem_AWBURST  = 2'b01;
    assign m07_axi_gmem_AWLOCK   = 2'b00;
    assign m07_axi_gmem_AWCACHE  = 4'b0011;
    assign m07_axi_gmem_AWPROT   = 3'b000;
    assign m07_axi_gmem_AWQOS    = 4'b0000;
    assign m07_axi_gmem_AWREGION = 4'b0000;
    assign m07_axi_gmem_ARBURST  = 2'b01;
    assign m07_axi_gmem_ARLOCK   = 2'b00;
    assign m07_axi_gmem_ARCACHE  = 4'b0011;
    assign m07_axi_gmem_ARPROT   = 3'b000;
    assign m07_axi_gmem_ARQOS    = 4'b0000;
    assign m07_axi_gmem_ARREGION = 4'b0000;

    assign m08_axi_gmem_AWID     = {C_M_AXI_GMEM_ID_WIDTH{1'b0}};
    assign m08_axi_gmem_AWBURST  = 2'b01;
    assign m08_axi_gmem_AWLOCK   = 2'b00;
    assign m08_axi_gmem_AWCACHE  = 4'b0011;
    assign m08_axi_gmem_AWPROT   = 3'b000;
    assign m08_axi_gmem_AWQOS    = 4'b0000;
    assign m08_axi_gmem_AWREGION = 4'b0000;
    assign m08_axi_gmem_ARBURST  = 2'b01;
    assign m08_axi_gmem_ARLOCK   = 2'b00;
    assign m08_axi_gmem_ARCACHE  = 4'b0011;
    assign m08_axi_gmem_ARPROT   = 3'b000;
    assign m08_axi_gmem_ARQOS    = 4'b0000;
    assign m08_axi_gmem_ARREGION = 4'b0000;

    assign m09_axi_gmem_AWID     = {C_M_AXI_GMEM_ID_WIDTH{1'b0}};
    assign m09_axi_gmem_AWBURST  = 2'b01;
    assign m09_axi_gmem_AWLOCK   = 2'b00;
    assign m09_axi_gmem_AWCACHE  = 4'b0011;
    assign m09_axi_gmem_AWPROT   = 3'b000;
    assign m09_axi_gmem_AWQOS    = 4'b0000;
    assign m09_axi_gmem_AWREGION = 4'b0000;
    assign m09_axi_gmem_ARBURST  = 2'b01;
    assign m09_axi_gmem_ARLOCK   = 2'b00;
    assign m09_axi_gmem_ARCACHE  = 4'b0011;
    assign m09_axi_gmem_ARPROT   = 3'b000;
    assign m09_axi_gmem_ARQOS    = 4'b0000;
    assign m09_axi_gmem_ARREGION = 4'b0000;

    assign m10_axi_gmem_AWID     = {C_M_AXI_GMEM_ID_WIDTH{1'b0}};
    assign m10_axi_gmem_AWBURST  = 2'b01;
    assign m10_axi_gmem_AWLOCK   = 2'b00;
    assign m10_axi_gmem_AWCACHE  = 4'b0011;
    assign m10_axi_gmem_AWPROT   = 3'b000;
    assign m10_axi_gmem_AWQOS    = 4'b0000;
    assign m10_axi_gmem_AWREGION = 4'b0000;
    assign m10_axi_gmem_ARBURST  = 2'b01;
    assign m10_axi_gmem_ARLOCK   = 2'b00;
    assign m10_axi_gmem_ARCACHE  = 4'b0011;
    assign m10_axi_gmem_ARPROT   = 3'b000;
    assign m10_axi_gmem_ARQOS    = 4'b0000;
    assign m10_axi_gmem_ARREGION = 4'b0000;

    assign m11_axi_gmem_AWID     = {C_M_AXI_GMEM_ID_WIDTH{1'b0}};
    assign m11_axi_gmem_AWBURST  = 2'b01;
    assign m11_axi_gmem_AWLOCK   = 2'b00;
    assign m11_axi_gmem_AWCACHE  = 4'b0011;
    assign m11_axi_gmem_AWPROT   = 3'b000;
    assign m11_axi_gmem_AWQOS    = 4'b0000;
    assign m11_axi_gmem_AWREGION = 4'b0000;
    assign m11_axi_gmem_ARBURST  = 2'b01;
    assign m11_axi_gmem_ARLOCK   = 2'b00;
    assign m11_axi_gmem_ARCACHE  = 4'b0011;
    assign m11_axi_gmem_ARPROT   = 3'b000;
    assign m11_axi_gmem_ARQOS    = 4'b0000;
    assign m11_axi_gmem_ARREGION = 4'b0000;

    assign m12_axi_gmem_AWID     = {C_M_AXI_GMEM_ID_WIDTH{1'b0}};
    assign m12_axi_gmem_AWBURST  = 2'b01;
    assign m12_axi_gmem_AWLOCK   = 2'b00;
    assign m12_axi_gmem_AWCACHE  = 4'b0011;
    assign m12_axi_gmem_AWPROT   = 3'b000;
    assign m12_axi_gmem_AWQOS    = 4'b0000;
    assign m12_axi_gmem_AWREGION = 4'b0000;
    assign m12_axi_gmem_ARBURST  = 2'b01;
    assign m12_axi_gmem_ARLOCK   = 2'b00;
    assign m12_axi_gmem_ARCACHE  = 4'b0011;
    assign m12_axi_gmem_ARPROT   = 3'b000;
    assign m12_axi_gmem_ARQOS    = 4'b0000;
    assign m12_axi_gmem_ARREGION = 4'b0000;

    assign m13_axi_gmem_AWID     = {C_M_AXI_GMEM_ID_WIDTH{1'b0}};
    assign m13_axi_gmem_AWBURST  = 2'b01;
    assign m13_axi_gmem_AWLOCK   = 2'b00;
    assign m13_axi_gmem_AWCACHE  = 4'b0011;
    assign m13_axi_gmem_AWPROT   = 3'b000;
    assign m13_axi_gmem_AWQOS    = 4'b0000;
    assign m13_axi_gmem_AWREGION = 4'b0000;
    assign m13_axi_gmem_ARBURST  = 2'b01;
    assign m13_axi_gmem_ARLOCK   = 2'b00;
    assign m13_axi_gmem_ARCACHE  = 4'b0011;
    assign m13_axi_gmem_ARPROT   = 3'b000;
    assign m13_axi_gmem_ARQOS    = 4'b0000;
    assign m13_axi_gmem_ARREGION = 4'b0000;

    assign m14_axi_gmem_AWID     = {C_M_AXI_GMEM_ID_WIDTH{1'b0}};
    assign m14_axi_gmem_AWBURST  = 2'b01;
    assign m14_axi_gmem_AWLOCK   = 2'b00;
    assign m14_axi_gmem_AWCACHE  = 4'b0011;
    assign m14_axi_gmem_AWPROT   = 3'b000;
    assign m14_axi_gmem_AWQOS    = 4'b0000;
    assign m14_axi_gmem_AWREGION = 4'b0000;
    assign m14_axi_gmem_ARBURST  = 2'b01;
    assign m14_axi_gmem_ARLOCK   = 2'b00;
    assign m14_axi_gmem_ARCACHE  = 4'b0011;
    assign m14_axi_gmem_ARPROT   = 3'b000;
    assign m14_axi_gmem_ARQOS    = 4'b0000;
    assign m14_axi_gmem_ARREGION = 4'b0000;

    assign m15_axi_gmem_AWID     = {C_M_AXI_GMEM_ID_WIDTH{1'b0}};
    assign m15_axi_gmem_AWBURST  = 2'b01;
    assign m15_axi_gmem_AWLOCK   = 2'b00;
    assign m15_axi_gmem_AWCACHE  = 4'b0011;
    assign m15_axi_gmem_AWPROT   = 3'b000;
    assign m15_axi_gmem_AWQOS    = 4'b0000;
    assign m15_axi_gmem_AWREGION = 4'b0000;
    assign m15_axi_gmem_ARBURST  = 2'b01;
    assign m15_axi_gmem_ARLOCK   = 2'b00;
    assign m15_axi_gmem_ARCACHE  = 4'b0011;
    assign m15_axi_gmem_ARPROT   = 3'b000;
    assign m15_axi_gmem_ARQOS    = 4'b0000;
    assign m15_axi_gmem_ARREGION = 4'b0000;

    assign m16_axi_gmem_AWID     = {C_M_AXI_GMEM_ID_WIDTH{1'b0}};
    assign m16_axi_gmem_AWBURST  = 2'b01;
    assign m16_axi_gmem_AWLOCK   = 2'b00;
    assign m16_axi_gmem_AWCACHE  = 4'b0011;
    assign m16_axi_gmem_AWPROT   = 3'b000;
    assign m16_axi_gmem_AWQOS    = 4'b0000;
    assign m16_axi_gmem_AWREGION = 4'b0000;
    assign m16_axi_gmem_ARBURST  = 2'b01;
    assign m16_axi_gmem_ARLOCK   = 2'b00;
    assign m16_axi_gmem_ARCACHE  = 4'b0011;
    assign m16_axi_gmem_ARPROT   = 3'b000;
    assign m16_axi_gmem_ARQOS    = 4'b0000;
    assign m16_axi_gmem_ARREGION = 4'b0000;

    assign m17_axi_gmem_AWID     = {C_M_AXI_GMEM_ID_WIDTH{1'b0}};
    assign m17_axi_gmem_AWBURST  = 2'b01;
    assign m17_axi_gmem_AWLOCK   = 2'b00;
    assign m17_axi_gmem_AWCACHE  = 4'b0011;
    assign m17_axi_gmem_AWPROT   = 3'b000;
    assign m17_axi_gmem_AWQOS    = 4'b0000;
    assign m17_axi_gmem_AWREGION = 4'b0000;
    assign m17_axi_gmem_ARBURST  = 2'b01;
    assign m17_axi_gmem_ARLOCK   = 2'b00;
    assign m17_axi_gmem_ARCACHE  = 4'b0011;
    assign m17_axi_gmem_ARPROT   = 3'b000;
    assign m17_axi_gmem_ARQOS    = 4'b0000;
    assign m17_axi_gmem_ARREGION = 4'b0000;

    assign m18_axi_gmem_AWID     = {C_M_AXI_GMEM_ID_WIDTH{1'b0}};
    assign m18_axi_gmem_AWBURST  = 2'b01;
    assign m18_axi_gmem_AWLOCK   = 2'b00;
    assign m18_axi_gmem_AWCACHE  = 4'b0011;
    assign m18_axi_gmem_AWPROT   = 3'b000;
    assign m18_axi_gmem_AWQOS    = 4'b0000;
    assign m18_axi_gmem_AWREGION = 4'b0000;
    assign m18_axi_gmem_ARBURST  = 2'b01;
    assign m18_axi_gmem_ARLOCK   = 2'b00;
    assign m18_axi_gmem_ARCACHE  = 4'b0011;
    assign m18_axi_gmem_ARPROT   = 3'b000;
    assign m18_axi_gmem_ARQOS    = 4'b0000;
    assign m18_axi_gmem_ARREGION = 4'b0000;

    assign m19_axi_gmem_AWID     = {C_M_AXI_GMEM_ID_WIDTH{1'b0}};
    assign m19_axi_gmem_AWBURST  = 2'b01;
    assign m19_axi_gmem_AWLOCK   = 2'b00;
    assign m19_axi_gmem_AWCACHE  = 4'b0011;
    assign m19_axi_gmem_AWPROT   = 3'b000;
    assign m19_axi_gmem_AWQOS    = 4'b0000;
    assign m19_axi_gmem_AWREGION = 4'b0000;
    assign m19_axi_gmem_ARBURST  = 2'b01;
    assign m19_axi_gmem_ARLOCK   = 2'b00;
    assign m19_axi_gmem_ARCACHE  = 4'b0011;
    assign m19_axi_gmem_ARPROT   = 3'b000;
    assign m19_axi_gmem_ARQOS    = 4'b0000;
    assign m19_axi_gmem_ARREGION = 4'b0000;

    assign m20_axi_gmem_AWID     = {C_M_AXI_GMEM_ID_WIDTH{1'b0}};
    assign m20_axi_gmem_AWBURST  = 2'b01;
    assign m20_axi_gmem_AWLOCK   = 2'b00;
    assign m20_axi_gmem_AWCACHE  = 4'b0011;
    assign m20_axi_gmem_AWPROT   = 3'b000;
    assign m20_axi_gmem_AWQOS    = 4'b0000;
    assign m20_axi_gmem_AWREGION = 4'b0000;
    assign m20_axi_gmem_ARBURST  = 2'b01;
    assign m20_axi_gmem_ARLOCK   = 2'b00;
    assign m20_axi_gmem_ARCACHE  = 4'b0011;
    assign m20_axi_gmem_ARPROT   = 3'b000;
    assign m20_axi_gmem_ARQOS    = 4'b0000;
    assign m20_axi_gmem_ARREGION = 4'b0000;

    assign m21_axi_gmem_AWID     = {C_M_AXI_GMEM_ID_WIDTH{1'b0}};
    assign m21_axi_gmem_AWBURST  = 2'b01;
    assign m21_axi_gmem_AWLOCK   = 2'b00;
    assign m21_axi_gmem_AWCACHE  = 4'b0011;
    assign m21_axi_gmem_AWPROT   = 3'b000;
    assign m21_axi_gmem_AWQOS    = 4'b0000;
    assign m21_axi_gmem_AWREGION = 4'b0000;
    assign m21_axi_gmem_ARBURST  = 2'b01;
    assign m21_axi_gmem_ARLOCK   = 2'b00;
    assign m21_axi_gmem_ARCACHE  = 4'b0011;
    assign m21_axi_gmem_ARPROT   = 3'b000;
    assign m21_axi_gmem_ARQOS    = 4'b0000;
    assign m21_axi_gmem_ARREGION = 4'b0000;

    assign m22_axi_gmem_AWID     = {C_M_AXI_GMEM_ID_WIDTH{1'b0}};
    assign m22_axi_gmem_AWBURST  = 2'b01;
    assign m22_axi_gmem_AWLOCK   = 2'b00;
    assign m22_axi_gmem_AWCACHE  = 4'b0011;
    assign m22_axi_gmem_AWPROT   = 3'b000;
    assign m22_axi_gmem_AWQOS    = 4'b0000;
    assign m22_axi_gmem_AWREGION = 4'b0000;
    assign m22_axi_gmem_ARBURST  = 2'b01;
    assign m22_axi_gmem_ARLOCK   = 2'b00;
    assign m22_axi_gmem_ARCACHE  = 4'b0011;
    assign m22_axi_gmem_ARPROT   = 3'b000;
    assign m22_axi_gmem_ARQOS    = 4'b0000;
    assign m22_axi_gmem_ARREGION = 4'b0000;

    assign m23_axi_gmem_AWID     = {C_M_AXI_GMEM_ID_WIDTH{1'b0}};
    assign m23_axi_gmem_AWBURST  = 2'b01;
    assign m23_axi_gmem_AWLOCK   = 2'b00;
    assign m23_axi_gmem_AWCACHE  = 4'b0011;
    assign m23_axi_gmem_AWPROT   = 3'b000;
    assign m23_axi_gmem_AWQOS    = 4'b0000;
    assign m23_axi_gmem_AWREGION = 4'b0000;
    assign m23_axi_gmem_ARBURST  = 2'b01;
    assign m23_axi_gmem_ARLOCK   = 2'b00;
    assign m23_axi_gmem_ARCACHE  = 4'b0011;
    assign m23_axi_gmem_ARPROT   = 3'b000;
    assign m23_axi_gmem_ARQOS    = 4'b0000;
    assign m23_axi_gmem_ARREGION = 4'b0000;

    assign m24_axi_gmem_AWID     = {C_M_AXI_GMEM_ID_WIDTH{1'b0}};
    assign m24_axi_gmem_AWBURST  = 2'b01;
    assign m24_axi_gmem_AWLOCK   = 2'b00;
    assign m24_axi_gmem_AWCACHE  = 4'b0011;
    assign m24_axi_gmem_AWPROT   = 3'b000;
    assign m24_axi_gmem_AWQOS    = 4'b0000;
    assign m24_axi_gmem_AWREGION = 4'b0000;
    assign m24_axi_gmem_ARBURST  = 2'b01;
    assign m24_axi_gmem_ARLOCK   = 2'b00;
    assign m24_axi_gmem_ARCACHE  = 4'b0011;
    assign m24_axi_gmem_ARPROT   = 3'b000;
    assign m24_axi_gmem_ARQOS    = 4'b0000;
    assign m24_axi_gmem_ARREGION = 4'b0000;

    assign m25_axi_gmem_AWID     = {C_M_AXI_GMEM_ID_WIDTH{1'b0}};
    assign m25_axi_gmem_AWBURST  = 2'b01;
    assign m25_axi_gmem_AWLOCK   = 2'b00;
    assign m25_axi_gmem_AWCACHE  = 4'b0011;
    assign m25_axi_gmem_AWPROT   = 3'b000;
    assign m25_axi_gmem_AWQOS    = 4'b0000;
    assign m25_axi_gmem_AWREGION = 4'b0000;
    assign m25_axi_gmem_ARBURST  = 2'b01;
    assign m25_axi_gmem_ARLOCK   = 2'b00;
    assign m25_axi_gmem_ARCACHE  = 4'b0011;
    assign m25_axi_gmem_ARPROT   = 3'b000;
    assign m25_axi_gmem_ARQOS    = 4'b0000;
    assign m25_axi_gmem_ARREGION = 4'b0000;

    assign m26_axi_gmem_AWID     = {C_M_AXI_GMEM_ID_WIDTH{1'b0}};
    assign m26_axi_gmem_AWBURST  = 2'b01;
    assign m26_axi_gmem_AWLOCK   = 2'b00;
    assign m26_axi_gmem_AWCACHE  = 4'b0011;
    assign m26_axi_gmem_AWPROT   = 3'b000;
    assign m26_axi_gmem_AWQOS    = 4'b0000;
    assign m26_axi_gmem_AWREGION = 4'b0000;
    assign m26_axi_gmem_ARBURST  = 2'b01;
    assign m26_axi_gmem_ARLOCK   = 2'b00;
    assign m26_axi_gmem_ARCACHE  = 4'b0011;
    assign m26_axi_gmem_ARPROT   = 3'b000;
    assign m26_axi_gmem_ARQOS    = 4'b0000;
    assign m26_axi_gmem_ARREGION = 4'b0000;

    assign m27_axi_gmem_AWID     = {C_M_AXI_GMEM_ID_WIDTH{1'b0}};
    assign m27_axi_gmem_AWBURST  = 2'b01;
    assign m27_axi_gmem_AWLOCK   = 2'b00;
    assign m27_axi_gmem_AWCACHE  = 4'b0011;
    assign m27_axi_gmem_AWPROT   = 3'b000;
    assign m27_axi_gmem_AWQOS    = 4'b0000;
    assign m27_axi_gmem_AWREGION = 4'b0000;
    assign m27_axi_gmem_ARBURST  = 2'b01;
    assign m27_axi_gmem_ARLOCK   = 2'b00;
    assign m27_axi_gmem_ARCACHE  = 4'b0011;
    assign m27_axi_gmem_ARPROT   = 3'b000;
    assign m27_axi_gmem_ARQOS    = 4'b0000;
    assign m27_axi_gmem_ARREGION = 4'b0000;

    assign m28_axi_gmem_AWID     = {C_M_AXI_GMEM_ID_WIDTH{1'b0}};
    assign m28_axi_gmem_AWBURST  = 2'b01;
    assign m28_axi_gmem_AWLOCK   = 2'b00;
    assign m28_axi_gmem_AWCACHE  = 4'b0011;
    assign m28_axi_gmem_AWPROT   = 3'b000;
    assign m28_axi_gmem_AWQOS    = 4'b0000;
    assign m28_axi_gmem_AWREGION = 4'b0000;
    assign m28_axi_gmem_ARBURST  = 2'b01;
    assign m28_axi_gmem_ARLOCK   = 2'b00;
    assign m28_axi_gmem_ARCACHE  = 4'b0011;
    assign m28_axi_gmem_ARPROT   = 3'b000;
    assign m28_axi_gmem_ARQOS    = 4'b0000;
    assign m28_axi_gmem_ARREGION = 4'b0000;

    assign m29_axi_gmem_AWID     = {C_M_AXI_GMEM_ID_WIDTH{1'b0}};
    assign m29_axi_gmem_AWBURST  = 2'b01;
    assign m29_axi_gmem_AWLOCK   = 2'b00;
    assign m29_axi_gmem_AWCACHE  = 4'b0011;
    assign m29_axi_gmem_AWPROT   = 3'b000;
    assign m29_axi_gmem_AWQOS    = 4'b0000;
    assign m29_axi_gmem_AWREGION = 4'b0000;
    assign m29_axi_gmem_ARBURST  = 2'b01;
    assign m29_axi_gmem_ARLOCK   = 2'b00;
    assign m29_axi_gmem_ARCACHE  = 4'b0011;
    assign m29_axi_gmem_ARPROT   = 3'b000;
    assign m29_axi_gmem_ARQOS    = 4'b0000;
    assign m29_axi_gmem_ARREGION = 4'b0000;

    assign m30_axi_gmem_AWID     = {C_M_AXI_GMEM_ID_WIDTH{1'b0}};
    assign m30_axi_gmem_AWBURST  = 2'b01;
    assign m30_axi_gmem_AWLOCK   = 2'b00;
    assign m30_axi_gmem_AWCACHE  = 4'b0011;
    assign m30_axi_gmem_AWPROT   = 3'b000;
    assign m30_axi_gmem_AWQOS    = 4'b0000;
    assign m30_axi_gmem_AWREGION = 4'b0000;
    assign m30_axi_gmem_ARBURST  = 2'b01;
    assign m30_axi_gmem_ARLOCK   = 2'b00;
    assign m30_axi_gmem_ARCACHE  = 4'b0011;
    assign m30_axi_gmem_ARPROT   = 3'b000;
    assign m30_axi_gmem_ARQOS    = 4'b0000;
    assign m30_axi_gmem_ARREGION = 4'b0000;

    assign m31_axi_gmem_AWID     = {C_M_AXI_GMEM_ID_WIDTH{1'b0}};
    assign m31_axi_gmem_AWBURST  = 2'b01;
    assign m31_axi_gmem_AWLOCK   = 2'b00;
    assign m31_axi_gmem_AWCACHE  = 4'b0011;
    assign m31_axi_gmem_AWPROT   = 3'b000;
    assign m31_axi_gmem_AWQOS    = 4'b0000;
    assign m31_axi_gmem_AWREGION = 4'b0000;
    assign m31_axi_gmem_ARBURST  = 2'b01;
    assign m31_axi_gmem_ARLOCK   = 2'b00;
    assign m31_axi_gmem_ARCACHE  = 4'b0011;
    assign m31_axi_gmem_ARPROT   = 3'b000;
    assign m31_axi_gmem_ARQOS    = 4'b0000;
    assign m31_axi_gmem_ARREGION = 4'b0000;

    // Register and invert reset signal for better timing.
    always @(posedge ap_clk) begin
        areset <= ~ap_rst_n;
    end

    // create pulse when ap_start transitions to 1
    always @(posedge ap_clk) begin
        begin
            ap_start_r <= ap_start;
        end
    end

    assign ap_start_pulse = ap_start & ~ap_start_r;

    // ap_idle is asserted when done is asserted, it is de-asserted when ap_start_pulse 
    // is asserted
    always @(posedge ap_clk) begin
        if (areset | dev_reset) begin
            ap_idle <= 1'b1;
        end
        else begin
            ap_idle <= ap_done        ? 1'b1 :
            ap_start_pulse ? 1'b0 :
            ap_idle;
        end
    end

    assign ap_ready = ap_done;

    // AXI4-Lite slave
    
    krnl_tsp_rtl_control_s_axi #(
    .C_S_AXI_ADDR_WIDTH( C_S_AXI_CONTROL_ADDR_WIDTH ),
    .C_S_AXI_DATA_WIDTH( C_S_AXI_CONTROL_DATA_WIDTH )
    )
    inst_krnl_tsp_control_s_axi (
        .AWVALID   ( s_axi_control_AWVALID         ) ,
        .AWREADY   ( s_axi_control_AWREADY         ) ,
        .AWADDR    ( s_axi_control_AWADDR          ) ,
        .WVALID    ( s_axi_control_WVALID          ) ,
        .WREADY    ( s_axi_control_WREADY          ) ,
        .WDATA     ( s_axi_control_WDATA           ) ,
        .WSTRB     ( s_axi_control_WSTRB           ) ,
        .ARVALID   ( s_axi_control_ARVALID         ) ,
        .ARREADY   ( s_axi_control_ARREADY         ) ,
        .ARADDR    ( s_axi_control_ARADDR          ) ,
        .RVALID    ( s_axi_control_RVALID          ) ,
        .RREADY    ( s_axi_control_RREADY          ) ,
        .RDATA     ( s_axi_control_RDATA           ) ,
        .RRESP     ( s_axi_control_RRESP           ) ,
        .BVALID    ( s_axi_control_BVALID          ) ,
        .BREADY    ( s_axi_control_BREADY          ) ,
        .BRESP     ( s_axi_control_BRESP           ) ,
        .ACLK      ( ap_clk                        ) ,
        .ARESET    ( areset | dev_reset            ) ,
        .ACLK_EN   ( 1'b1                          ) ,
        .ap_start  ( ap_start                      ) ,
        .interrupt ( interrupt                     ) ,
        .ap_ready  ( ap_ready                      ) ,
        .ap_done   ( ap_done                       ) ,
        .ap_idle   ( ap_idle                       ) ,
        // User signals
        .file_size      ( file_size  ) ,
        .load_filesize  ( ctrl_load_filesize ) ,
        .start_address  ( start_addr ) ,
        .load_address   ( ctrl_load_address  ) ,
        .next_filesize  ( fm_next_filesize ) ,
        .next_address   ( fm_next_address ) ,
        .overlap        ( fm_overlap ) ,
        //.load_done      ( fm_done ) ,
        .load_done      ( &rd_channel_idle ) ,
        .dev_reset      ( dev_reset ),
        .dev_continue   ( dev_continue ) ,
        .dev_bytemode   ( dev_bytemode ) ,
        .dev_done       ( dev_done ) ,
        .dev_start      ( dev_start ) ,
        .dev_load_text  ( dev_load_text ) ,
        .key            ( ikey ) ,
        .key_we         ( ikey_wren ),
        .rden           ( result_rden ) ,
        .keylen         ( key_len ) ,
        .result         ( { result_valid, result_data } ),
        .bitstream_rden ( bitstream_rden           ),
        .bitsream       ( bitstream),
        .matchcount     ( match_count ),
        .matchcount_vld ( match_count_vld ),
        .bash_offset    ( fm_bash_offset   ) ,
        .bash_code      ( fm_bashcount     ) ,
        .bash_update    ( fm_bashupdate )
    );

    file_manager file_manager_inst(
        .clk            ( ap_clk             ) ,
        .reset          ( areset | dev_reset ) ,
        .istart         ( dev_load_text      ) ,
        .iload          ( ctrl_load_filesize ) ,
        .iload_address  ( ctrl_load_address  ) ,
        .idone          ( rd_done            ) ,
        .start_address  ( start_addr         ) ,
        .file_size      ( file_size          ) ,
        .ostart         ( load_start         ) ,
        .oreset         ( rd_reset           ) ,
        .ready          ( fm_ready           ) ,
        .odone          ( fm_done            ) ,
        .ofilesize      ( fm_next_filesize   ) ,
        .onext_addr     ( fm_next_address    ) ,
        .bash_offset    ( fm_bash_offset     ) ,          
        .bash_count     ( fm_bashcount       ) ,
        .bash_update    ( fm_bashupdate      ) ,
        .overlap        ( fm_overlap         ) ,
        .oc0_addr       ( rd_addr[0]         ) ,
        .oc1_addr       ( rd_addr[1]         ) ,
        .oc2_addr       ( rd_addr[2]         ) ,
        .oc3_addr       ( rd_addr[3]         ) ,
        .oc4_addr       ( rd_addr[4]         ) ,
        .oc5_addr       ( rd_addr[5]         ) ,
        .oc6_addr       ( rd_addr[6]         ) ,
        .oc7_addr       ( rd_addr[7]         ) ,
        .oc8_addr       ( rd_addr[8]         ) ,
        .oc9_addr       ( rd_addr[9]         ) ,
        .oc10_addr      ( rd_addr[10]        ) ,
        .oc11_addr      ( rd_addr[11]        ) ,
        .oc12_addr      ( rd_addr[12]        ) ,
        .oc13_addr      ( rd_addr[13]        ) ,
        .oc14_addr      ( rd_addr[14]        ) ,
        .oc15_addr      ( rd_addr[15]        ) ,
        .oc16_addr      ( rd_addr[16]        ) ,
        .oc17_addr      ( rd_addr[17]        ) ,
        .oc18_addr      ( rd_addr[18]        ) ,
        .oc19_addr      ( rd_addr[19]        ) ,
        .oc20_addr      ( rd_addr[20]        ) ,
        .oc21_addr      ( rd_addr[21]        ) ,
        .oc22_addr      ( rd_addr[22]        ) ,
        .oc23_addr      ( rd_addr[23]        ) ,
        .oc24_addr      ( rd_addr[24]        ) ,
        .oc25_addr      ( rd_addr[25]        ) ,
        .oc26_addr      ( rd_addr[26]        ) ,
        .oc27_addr      ( rd_addr[27]        ) ,
        .oc28_addr      ( rd_addr[28]        ) ,
        .oc29_addr      ( rd_addr[29]        ) ,
        .oc30_addr      ( rd_addr[30]        ) ,
        .oc31_addr      ( rd_addr[31]        ) ,
        .oc0_rdlen      ( rd_length[0]       ) ,
        .oc1_rdlen      ( rd_length[1]       ) ,
        .oc2_rdlen      ( rd_length[2]       ) ,
        .oc3_rdlen      ( rd_length[3]       ) ,
        .oc4_rdlen      ( rd_length[4]       ) ,
        .oc5_rdlen      ( rd_length[5]       ) ,
        .oc6_rdlen      ( rd_length[6]       ) ,
        .oc7_rdlen      ( rd_length[7]       ) ,
        .oc8_rdlen      ( rd_length[8]       ) ,
        .oc9_rdlen      ( rd_length[9]       ) ,
        .oc10_rdlen     ( rd_length[10]      ) ,
        .oc11_rdlen     ( rd_length[11]      ) ,
        .oc12_rdlen     ( rd_length[12]      ) ,
        .oc13_rdlen     ( rd_length[13]      ) ,
        .oc14_rdlen     ( rd_length[14]      ) ,
        .oc15_rdlen     ( rd_length[15]      ) ,
        .oc16_rdlen     ( rd_length[16]      ) ,
        .oc17_rdlen     ( rd_length[17]      ) ,
        .oc18_rdlen     ( rd_length[18]      ) ,
        .oc19_rdlen     ( rd_length[19]      ) ,
        .oc20_rdlen     ( rd_length[20]      ) ,
        .oc21_rdlen     ( rd_length[21]      ) ,
        .oc22_rdlen     ( rd_length[22]      ) ,
        .oc23_rdlen     ( rd_length[23]      ) ,
        .oc24_rdlen     ( rd_length[24]      ) ,
        .oc25_rdlen     ( rd_length[25]      ) ,
        .oc26_rdlen     ( rd_length[26]      ) ,
        .oc27_rdlen     ( rd_length[27]      ) ,
        .oc28_rdlen     ( rd_length[28]      ) ,
        .oc29_rdlen     ( rd_length[29]      ) ,
        .oc30_rdlen     ( rd_length[30]      ) ,
        .oc31_rdlen     ( rd_length[31]      )
    );

    krnl_rtl_read_axi #(
    .C_ADDR_WIDTH     ( C_M_AXI_GMEM_ADDR_WIDTH ) ,
    .C_DATA_WIDTH     ( C_M_AXI_GMEM_DATA_WIDTH ) ,
    .C_LENGTH_WIDTH   ( LP_LENGTH_WIDTH         ) ,
    .C_BURST_LEN      ( LP_AXI_BURST_LEN        ) ,
    .C_LOG_BURST_LEN  ( LP_LOG_BURST_LEN        ) ,
    .C_MAX_OUTSTANDING( LP_RD_MAX_OUTSTANDING   )
    )
    axi_read_master_inst00(
        // System signals
        .aclk         ( ap_clk ) , // input
        .areset       ( areset | dev_load_text | dev_continue | dev_reset) , // input
        // Control signals 
        .dev_start    ( fm_done    ) ,
        .load_done    ( fm_done    ) ,
        .ctrl_start   ( load_start[0]) , // input
        .ctrl_done    ( rd_done[0]   ) , // output
        .ctrl_offset  ( rd_addr[0]   ) , // input [C_ADDR_WIDTH-1:0]
        .ctrl_length  ( rd_length[0] ) , // input [C_LENGTH_WIDTH-1:0]
        // AXI4 master interface                             
        .arvalid      ( m00_axi_gmem_ARVALID ) , // output
        .arready      ( m00_axi_gmem_ARREADY ) , // input
        .araddr       ( m00_axi_gmem_ARADDR  ) , // output [C_ADDR_WIDTH-1:0]
        .arid         ( m00_axi_gmem_ARID    ) , // output
        .arlen        ( m00_axi_gmem_ARLEN   ) , // output
        .arsize       ( m00_axi_gmem_ARSIZE  ) , // output [2:0]
        .rvalid       ( m00_axi_gmem_RVALID  ) , // input
        .rready       ( m00_axi_gmem_RREADY  ) , // output
        .rdata        ( m00_axi_gmem_RDATA   ) , // input [C_DATA_WIDTH - 1:0]
        .rlast        ( m00_axi_gmem_RLAST   ) , // input
        .rid          ( m00_axi_gmem_RID     ) , // input
        .rresp        ( m00_axi_gmem_RRESP   ) , // input [1:0]
        // FIFO read signals
        .idle         ( rd_channel_idle[0]   ) ,  
        .odone        ( rd_done2[0]          ) ,
        .rd_en        ( rd_en[0]             ) , // input
        .rd_data      ( rd_data[0]           ) , // output [C_DATA_WIDTH - 1:0]
        .rd_tvalid_n  ( rd_tvalid_n[0]       ) ,// output
        .ocount       ( count0[7:0] ),
        .ostate       ( count1[7:0] )
    );

    krnl_rtl_read_axi #(
    .C_ADDR_WIDTH     ( C_M_AXI_GMEM_ADDR_WIDTH ) ,
    .C_DATA_WIDTH     ( C_M_AXI_GMEM_DATA_WIDTH ) ,
    .C_LENGTH_WIDTH   ( LP_LENGTH_WIDTH         ) ,
    .C_BURST_LEN      ( LP_AXI_BURST_LEN        ) ,
    .C_LOG_BURST_LEN  ( LP_LOG_BURST_LEN        ) ,
    .C_MAX_OUTSTANDING( LP_RD_MAX_OUTSTANDING   )
    )
    axi_read_master_inst01(
        // System signals
        .aclk         ( ap_clk ) , // input
        .areset       ( rd_reset | dev_load_text |  dev_continue | dev_reset ) , // input
        // Control signals 
        .dev_start    ( fm_done       ) ,
        .load_done    ( fm_done       ) ,
        .ctrl_start   ( load_start[1]   ) , // input
        .ctrl_done    ( rd_done[1]      ) , // output
        .ctrl_offset  ( rd_addr[1]      ) , // input [C_ADDR_WIDTH-1:0]
        .ctrl_length  ( rd_length[1]    ) , // input [C_LENGTH_WIDTH-1:0]
        // AXI4 master interface                             
        .arvalid      ( m01_axi_gmem_ARVALID ) , // output
        .arready      ( m01_axi_gmem_ARREADY ) , // input
        .araddr       ( m01_axi_gmem_ARADDR  ) , // output [C_ADDR_WIDTH-1:0]
        .arid         ( m01_axi_gmem_ARID    ) , // output
        .arlen        ( m01_axi_gmem_ARLEN   ) , // output
        .arsize       ( m01_axi_gmem_ARSIZE  ) , // output [2:0]
        .rvalid       ( m01_axi_gmem_RVALID  ) , // input
        .rready       ( m01_axi_gmem_RREADY  ) , // output
        .rdata        ( m01_axi_gmem_RDATA   ) , // input [C_DATA_WIDTH - 1:0]
        .rlast        ( m01_axi_gmem_RLAST   ) , // input
        .rid          ( m01_axi_gmem_RID     ) , // input
        .rresp        ( m01_axi_gmem_RRESP   ) , // input [1:0]
        // FIFO read signals
        .idle         ( rd_channel_idle[1]   ) ,
        .odone        ( rd_done2[1]          ) ,
        .rd_en        ( rd_en[1]             ) , // input
        .rd_data      ( rd_data[1]           ) , // output [C_DATA_WIDTH - 1:0]
        .rd_tvalid_n  ( rd_tvalid_n[1]       ) ,// output
        .ocount       ( count0[15:8] ),
        .ostate       ( count1[15:8] )
    );

    krnl_rtl_read_axi #(
    .C_ADDR_WIDTH     ( C_M_AXI_GMEM_ADDR_WIDTH ) ,
    .C_DATA_WIDTH     ( C_M_AXI_GMEM_DATA_WIDTH ) ,
    .C_LENGTH_WIDTH   ( LP_LENGTH_WIDTH         ) ,
    .C_BURST_LEN      ( LP_AXI_BURST_LEN        ) ,
    .C_LOG_BURST_LEN  ( LP_LOG_BURST_LEN        ) ,
    .C_MAX_OUTSTANDING( LP_RD_MAX_OUTSTANDING   )
    )
    axi_read_master_inst02(
        // System signals
        .aclk         ( ap_clk ) , // input
        .areset       ( rd_reset | dev_load_text |  dev_continue | dev_reset ) , // input
        // Control signals 
        .dev_start    ( fm_done       ) ,
        .load_done    ( fm_done       ) ,
        .ctrl_start   ( load_start[2]   ) , // input
        .ctrl_done    ( rd_done[2]      ) , // output
        .ctrl_offset  ( rd_addr[2]      ) , // input [C_ADDR_WIDTH-1:0]
        .ctrl_length  ( rd_length[2]    ) , // input [C_LENGTH_WIDTH-1:0]
        // AXI4 master interface                             
        .arvalid      ( m02_axi_gmem_ARVALID ) , // output
        .arready      ( m02_axi_gmem_ARREADY ) , // input
        .araddr       ( m02_axi_gmem_ARADDR  ) , // output [C_ADDR_WIDTH-1:0]
        .arid         ( m02_axi_gmem_ARID    ) , // output
        .arlen        ( m02_axi_gmem_ARLEN   ) , // output
        .arsize       ( m02_axi_gmem_ARSIZE  ) , // output [2:0]
        .rvalid       ( m02_axi_gmem_RVALID  ) , // input
        .rready       ( m02_axi_gmem_RREADY  ) , // output
        .rdata        ( m02_axi_gmem_RDATA   ) , // input [C_DATA_WIDTH - 1:0]
        .rlast        ( m02_axi_gmem_RLAST   ) , // input
        .rid          ( m02_axi_gmem_RID     ) , // input
        .rresp        ( m02_axi_gmem_RRESP   ) , // input [1:0]
        // FIFO read signals
        .idle         ( rd_channel_idle[2]   ) ,
        .odone        ( rd_done2[2]          ) ,
        .rd_en        ( rd_en[2]             ) , // input
        .rd_data      ( rd_data[2]           ) , // output [C_DATA_WIDTH - 1:0]
        .rd_tvalid_n  ( rd_tvalid_n[2]       ) // output
    );

    krnl_rtl_read_axi #(
    .C_ADDR_WIDTH     ( C_M_AXI_GMEM_ADDR_WIDTH ) ,
    .C_DATA_WIDTH     ( C_M_AXI_GMEM_DATA_WIDTH ) ,
    .C_LENGTH_WIDTH   ( LP_LENGTH_WIDTH         ) ,
    .C_BURST_LEN      ( LP_AXI_BURST_LEN        ) ,
    .C_LOG_BURST_LEN  ( LP_LOG_BURST_LEN        ) ,
    .C_MAX_OUTSTANDING( LP_RD_MAX_OUTSTANDING   )
    )
    axi_read_master_inst03(
        // System signals
        .aclk         ( ap_clk ) , // input
        .areset       ( rd_reset | dev_load_text |  dev_continue | dev_reset ) , // input
        // Control signals 
        .dev_start    ( fm_done       ) ,
        .load_done    ( fm_done       ) ,
        .ctrl_start   ( load_start[3]   ) , // input
        .ctrl_done    ( rd_done[3]      ) , // output
        .ctrl_offset  ( rd_addr[3]      ) , // input [C_ADDR_WIDTH-1:0]
        .ctrl_length  ( rd_length[3]    ) , // input [C_LENGTH_WIDTH-1:0]
        // AXI4 master interface                             
        .arvalid      ( m03_axi_gmem_ARVALID ) , // output
        .arready      ( m03_axi_gmem_ARREADY ) , // input
        .araddr       ( m03_axi_gmem_ARADDR  ) , // output [C_ADDR_WIDTH-1:0]
        .arid         ( m03_axi_gmem_ARID    ) , // output
        .arlen        ( m03_axi_gmem_ARLEN   ) , // output
        .arsize       ( m03_axi_gmem_ARSIZE  ) , // output [2:0]
        .rvalid       ( m03_axi_gmem_RVALID  ) , // input
        .rready       ( m03_axi_gmem_RREADY  ) , // output
        .rdata        ( m03_axi_gmem_RDATA   ) , // input [C_DATA_WIDTH - 1:0]
        .rlast        ( m03_axi_gmem_RLAST   ) , // input
        .rid          ( m03_axi_gmem_RID     ) , // input
        .rresp        ( m03_axi_gmem_RRESP   ) , // input [1:0]
        // FIFO read signals
        .idle         ( rd_channel_idle[3]   ) ,
        .odone        ( rd_done2[3]          ) ,
        .rd_en        ( rd_en[3]             ) , // input
        .rd_data      ( rd_data[3]           ) , // output [C_DATA_WIDTH - 1:0]
        .rd_tvalid_n  ( rd_tvalid_n[3]       ) // output
    );

    krnl_rtl_read_axi #(
    .C_ADDR_WIDTH     ( C_M_AXI_GMEM_ADDR_WIDTH ) ,
    .C_DATA_WIDTH     ( C_M_AXI_GMEM_DATA_WIDTH ) ,
    .C_LENGTH_WIDTH   ( LP_LENGTH_WIDTH         ) ,
    .C_BURST_LEN      ( LP_AXI_BURST_LEN        ) ,
    .C_LOG_BURST_LEN  ( LP_LOG_BURST_LEN        ) ,
    .C_MAX_OUTSTANDING( LP_RD_MAX_OUTSTANDING   )
    )
    axi_read_master_inst04(
        // System signals
        .aclk         ( ap_clk ) , // input
        .areset       ( rd_reset | dev_load_text |  dev_continue | dev_reset ) , // input
        // Control signals 
        .dev_start    ( fm_done) ,
        .load_done    ( fm_done      ) ,
        .ctrl_start   ( load_start[4] ) , // input
        .ctrl_done    ( rd_done[4]      ) , // output
        .ctrl_offset  ( rd_addr[4]      ) , // input [C_ADDR_WIDTH-1:0]
        .ctrl_length  ( rd_length[4]    ) , // input [C_LENGTH_WIDTH-1:0]
        // AXI4 master interface                             
        .arvalid      ( m04_axi_gmem_ARVALID ) , // output
        .arready      ( m04_axi_gmem_ARREADY ) , // input
        .araddr       ( m04_axi_gmem_ARADDR  ) , // output [C_ADDR_WIDTH-1:0]
        .arid         ( m04_axi_gmem_ARID    ) , // output
        .arlen        ( m04_axi_gmem_ARLEN   ) , // output
        .arsize       ( m04_axi_gmem_ARSIZE  ) , // output [2:0]
        .rvalid       ( m04_axi_gmem_RVALID  ) , // input
        .rready       ( m04_axi_gmem_RREADY  ) , // output
        .rdata        ( m04_axi_gmem_RDATA   ) , // input [C_DATA_WIDTH - 1:0]
        .rlast        ( m04_axi_gmem_RLAST   ) , // input
        .rid          ( m04_axi_gmem_RID     ) , // input
        .rresp        ( m04_axi_gmem_RRESP   ) , // input [1:0]
        // FIFO read signals
        .idle         ( rd_channel_idle[4]   ) ,
        .odone        ( rd_done2[4]          ) ,
        .rd_en        ( rd_en[4]             ) , // input
        .rd_data      ( rd_data[4]           ) , // output [C_DATA_WIDTH - 1:0]
        .rd_tvalid_n  ( rd_tvalid_n[4]       ) // output
    );

    krnl_rtl_read_axi #(
    .C_ADDR_WIDTH     ( C_M_AXI_GMEM_ADDR_WIDTH ) ,
    .C_DATA_WIDTH     ( C_M_AXI_GMEM_DATA_WIDTH ) ,
    .C_LENGTH_WIDTH   ( LP_LENGTH_WIDTH         ) ,
    .C_BURST_LEN      ( LP_AXI_BURST_LEN        ) ,
    .C_LOG_BURST_LEN  ( LP_LOG_BURST_LEN        ) ,
    .C_MAX_OUTSTANDING( LP_RD_MAX_OUTSTANDING   )
    )
    axi_read_master_inst05(
        // System signals
        .aclk         ( ap_clk ) , // input
        .areset       ( rd_reset | dev_load_text |  dev_continue | dev_reset ) , // input
        // Control signals 
        .dev_start    ( fm_done) ,
        .load_done    ( fm_done      ) ,
        .ctrl_start   ( load_start[5] ) , // input
        .ctrl_done    ( rd_done[5]      ) , // output
        .ctrl_offset  ( rd_addr[5]      ) , // input [C_ADDR_WIDTH-1:0]
        .ctrl_length  ( rd_length[5]    ) , // input [C_LENGTH_WIDTH-1:0]
        // AXI4 master interface                             
        .arvalid      ( m05_axi_gmem_ARVALID ) , // output
        .arready      ( m05_axi_gmem_ARREADY ) , // input
        .araddr       ( m05_axi_gmem_ARADDR  ) , // output [C_ADDR_WIDTH-1:0]
        .arid         ( m05_axi_gmem_ARID    ) , // output
        .arlen        ( m05_axi_gmem_ARLEN   ) , // output
        .arsize       ( m05_axi_gmem_ARSIZE  ) , // output [2:0]
        .rvalid       ( m05_axi_gmem_RVALID  ) , // input
        .rready       ( m05_axi_gmem_RREADY  ) , // output
        .rdata        ( m05_axi_gmem_RDATA   ) , // input [C_DATA_WIDTH - 1:0]
        .rlast        ( m05_axi_gmem_RLAST   ) , // input
        .rid          ( m05_axi_gmem_RID     ) , // input
        .rresp        ( m05_axi_gmem_RRESP   ) , // input [1:0]
        // FIFO read signals
        .idle         ( rd_channel_idle[5]   ) ,
        .odone        ( rd_done2[5]          ) ,
        .rd_en        ( rd_en[5]             ) , // input
        .rd_data      ( rd_data[5]           ) , // output [C_DATA_WIDTH - 1:0]
        .rd_tvalid_n  ( rd_tvalid_n[5]       ) // output
    );

    krnl_rtl_read_axi #(
    .C_ADDR_WIDTH     ( C_M_AXI_GMEM_ADDR_WIDTH ) ,
    .C_DATA_WIDTH     ( C_M_AXI_GMEM_DATA_WIDTH ) ,
    .C_LENGTH_WIDTH   ( LP_LENGTH_WIDTH         ) ,
    .C_BURST_LEN      ( LP_AXI_BURST_LEN        ) ,
    .C_LOG_BURST_LEN  ( LP_LOG_BURST_LEN        ) ,
    .C_MAX_OUTSTANDING( LP_RD_MAX_OUTSTANDING   )
    )
    axi_read_master_inst06(
        // System signals
        .aclk         ( ap_clk ) , // input
        .areset       ( rd_reset | dev_load_text |  dev_continue | dev_reset ) , // input
        // Control signals 
        .dev_start    ( fm_done) ,
        .load_done    ( fm_done      ) ,
        .ctrl_start   ( load_start[6] ) , // input
        .ctrl_done    ( rd_done[6]      ) , // output
        .ctrl_offset  ( rd_addr[6]      ) , // input [C_ADDR_WIDTH-1:0]
        .ctrl_length  ( rd_length[6]    ) , // input [C_LENGTH_WIDTH-1:0]
        // AXI4 master interface                             
        .arvalid      ( m06_axi_gmem_ARVALID ) , // output
        .arready      ( m06_axi_gmem_ARREADY ) , // input
        .araddr       ( m06_axi_gmem_ARADDR  ) , // output [C_ADDR_WIDTH-1:0]
        .arid         ( m06_axi_gmem_ARID    ) , // output
        .arlen        ( m06_axi_gmem_ARLEN   ) , // output
        .arsize       ( m06_axi_gmem_ARSIZE  ) , // output [2:0]
        .rvalid       ( m06_axi_gmem_RVALID  ) , // input
        .rready       ( m06_axi_gmem_RREADY  ) , // output
        .rdata        ( m06_axi_gmem_RDATA   ) , // input [C_DATA_WIDTH - 1:0]
        .rlast        ( m06_axi_gmem_RLAST   ) , // input
        .rid          ( m06_axi_gmem_RID     ) , // input
        .rresp        ( m06_axi_gmem_RRESP   ) , // input [1:0]
        // FIFO read signals
        .idle         ( rd_channel_idle[6]   ) ,
        .odone        ( rd_done2[6]          ) ,
        .rd_en        ( rd_en[6]             ) , // input
        .rd_data      ( rd_data[6]           ) , // output [C_DATA_WIDTH - 1:0]
        .rd_tvalid_n  ( rd_tvalid_n[6]       ) // output
    );

    krnl_rtl_read_axi #(
    .C_ADDR_WIDTH     ( C_M_AXI_GMEM_ADDR_WIDTH ) ,
    .C_DATA_WIDTH     ( C_M_AXI_GMEM_DATA_WIDTH ) ,
    .C_LENGTH_WIDTH   ( LP_LENGTH_WIDTH         ) ,
    .C_BURST_LEN      ( LP_AXI_BURST_LEN        ) ,
    .C_LOG_BURST_LEN  ( LP_LOG_BURST_LEN        ) ,
    .C_MAX_OUTSTANDING( LP_RD_MAX_OUTSTANDING   )
    )
    axi_read_master_inst07(
        // System signals
        .aclk         ( ap_clk ) , // input
        .areset       ( rd_reset | dev_load_text |  dev_continue | dev_reset ) , // input
        // Control signals 
        .dev_start    ( fm_done) ,
        .load_done    ( fm_done      ) ,
        .ctrl_start   ( load_start[7] ) , // input
        .ctrl_done    ( rd_done[7]      ) , // output
        .ctrl_offset  ( rd_addr[7]      ) , // input [C_ADDR_WIDTH-1:0]
        .ctrl_length  ( rd_length[7]    ) , // input [C_LENGTH_WIDTH-1:0]
        // AXI4 master interface                             
        .arvalid      ( m07_axi_gmem_ARVALID ) , // output
        .arready      ( m07_axi_gmem_ARREADY ) , // input
        .araddr       ( m07_axi_gmem_ARADDR  ) , // output [C_ADDR_WIDTH-1:0]
        .arid         ( m07_axi_gmem_ARID    ) , // output
        .arlen        ( m07_axi_gmem_ARLEN   ) , // output
        .arsize       ( m07_axi_gmem_ARSIZE  ) , // output [2:0]
        .rvalid       ( m07_axi_gmem_RVALID  ) , // input
        .rready       ( m07_axi_gmem_RREADY  ) , // output
        .rdata        ( m07_axi_gmem_RDATA   ) , // input [C_DATA_WIDTH - 1:0]
        .rlast        ( m07_axi_gmem_RLAST   ) , // input
        .rid          ( m07_axi_gmem_RID     ) , // input
        .rresp        ( m07_axi_gmem_RRESP   ) , // input [1:0]
        // FIFO read signals
        .idle         ( rd_channel_idle[7]   ) ,
        .odone        ( rd_done2[7]          ) ,
        .rd_en        ( rd_en[7]             ) , // input
        .rd_data      ( rd_data[7]           ) , // output [C_DATA_WIDTH - 1:0]
        .rd_tvalid_n  ( rd_tvalid_n[7]       ) // output
    );

    krnl_rtl_read_axi #(
    .C_ADDR_WIDTH     ( C_M_AXI_GMEM_ADDR_WIDTH ) ,
    .C_DATA_WIDTH     ( C_M_AXI_GMEM_DATA_WIDTH ) ,
    .C_LENGTH_WIDTH   ( LP_LENGTH_WIDTH         ) ,
    .C_BURST_LEN      ( LP_AXI_BURST_LEN        ) ,
    .C_LOG_BURST_LEN  ( LP_LOG_BURST_LEN        ) ,
    .C_MAX_OUTSTANDING( LP_RD_MAX_OUTSTANDING   )
    )
    axi_read_master_inst08(
        // System signals
        .aclk         ( ap_clk ) , // input
        .areset       ( rd_reset | dev_load_text |  dev_continue | dev_reset ) , // input
        // Control signals 
        .dev_start    ( fm_done) ,
        .load_done    ( fm_done      ) ,
        .ctrl_start   ( load_start[8] ) , // input
        .ctrl_done    ( rd_done[8]      ) , // output
        .ctrl_offset  ( rd_addr[8]      ) , // input [C_ADDR_WIDTH-1:0]
        .ctrl_length  ( rd_length[8]    ) , // input [C_LENGTH_WIDTH-1:0]
        // AXI4 master interface                             
        .arvalid      ( m08_axi_gmem_ARVALID ) , // output
        .arready      ( m08_axi_gmem_ARREADY ) , // input
        .araddr       ( m08_axi_gmem_ARADDR  ) , // output [C_ADDR_WIDTH-1:0]
        .arid         ( m08_axi_gmem_ARID    ) , // output
        .arlen        ( m08_axi_gmem_ARLEN   ) , // output
        .arsize       ( m08_axi_gmem_ARSIZE  ) , // output [2:0]
        .rvalid       ( m08_axi_gmem_RVALID  ) , // input
        .rready       ( m08_axi_gmem_RREADY  ) , // output
        .rdata        ( m08_axi_gmem_RDATA   ) , // input [C_DATA_WIDTH - 1:0]
        .rlast        ( m08_axi_gmem_RLAST   ) , // input
        .rid          ( m08_axi_gmem_RID     ) , // input
        .rresp        ( m08_axi_gmem_RRESP   ) , // input [1:0]
        // FIFO read signals
        .idle         ( rd_channel_idle[8]   ) ,
        .odone        ( rd_done2[8]          ) ,
        .rd_en        ( rd_en[8]             ) , // input
        .rd_data      ( rd_data[8]           ) , // output [C_DATA_WIDTH - 1:0]
        .rd_tvalid_n  ( rd_tvalid_n[8]       ) // output
    );

    krnl_rtl_read_axi #(
    .C_ADDR_WIDTH     ( C_M_AXI_GMEM_ADDR_WIDTH ) ,
    .C_DATA_WIDTH     ( C_M_AXI_GMEM_DATA_WIDTH ) ,
    .C_LENGTH_WIDTH   ( LP_LENGTH_WIDTH         ) ,
    .C_BURST_LEN      ( LP_AXI_BURST_LEN        ) ,
    .C_LOG_BURST_LEN  ( LP_LOG_BURST_LEN        ) ,
    .C_MAX_OUTSTANDING( LP_RD_MAX_OUTSTANDING   )
    )
    axi_read_master_inst09(
        // System signals
        .aclk         ( ap_clk ) , // input
        .areset       ( rd_reset | dev_load_text |  dev_continue | dev_reset ) , // input
        // Control signals 
        .dev_start    ( fm_done) ,
        .load_done    ( fm_done      ) ,
        .ctrl_start   ( load_start[9] ) , // input
        .ctrl_done    ( rd_done[9]      ) , // output
        .ctrl_offset  ( rd_addr[9]      ) , // input [C_ADDR_WIDTH-1:0]
        .ctrl_length  ( rd_length[9]    ) , // input [C_LENGTH_WIDTH-1:0]
        // AXI4 master interface                             
        .arvalid      ( m09_axi_gmem_ARVALID ) , // output
        .arready      ( m09_axi_gmem_ARREADY ) , // input
        .araddr       ( m09_axi_gmem_ARADDR  ) , // output [C_ADDR_WIDTH-1:0]
        .arid         ( m09_axi_gmem_ARID    ) , // output
        .arlen        ( m09_axi_gmem_ARLEN   ) , // output
        .arsize       ( m09_axi_gmem_ARSIZE  ) , // output [2:0]
        .rvalid       ( m09_axi_gmem_RVALID  ) , // input
        .rready       ( m09_axi_gmem_RREADY  ) , // output
        .rdata        ( m09_axi_gmem_RDATA   ) , // input [C_DATA_WIDTH - 1:0]
        .rlast        ( m09_axi_gmem_RLAST   ) , // input
        .rid          ( m09_axi_gmem_RID     ) , // input
        .rresp        ( m09_axi_gmem_RRESP   ) , // input [1:0]
        // FIFO read signals
        .idle         ( rd_channel_idle[9]   ) ,
        .odone        ( rd_done2[9]          ) ,
        .rd_en        ( rd_en[9]             ) , // input
        .rd_data      ( rd_data[9]           ) , // output [C_DATA_WIDTH - 1:0]
        .rd_tvalid_n  ( rd_tvalid_n[9]       ) // output
    );

    krnl_rtl_read_axi #(
    .C_ADDR_WIDTH     ( C_M_AXI_GMEM_ADDR_WIDTH ) ,
    .C_DATA_WIDTH     ( C_M_AXI_GMEM_DATA_WIDTH ) ,
    .C_LENGTH_WIDTH   ( LP_LENGTH_WIDTH         ) ,
    .C_BURST_LEN      ( LP_AXI_BURST_LEN        ) ,
    .C_LOG_BURST_LEN  ( LP_LOG_BURST_LEN        ) ,
    .C_MAX_OUTSTANDING( LP_RD_MAX_OUTSTANDING   )
    )
    axi_read_master_inst10(
        // System signals
        .aclk         ( ap_clk ) , // input
        .areset       ( rd_reset | dev_load_text |  dev_continue | dev_reset ) , // input
        // Control signals 
        .dev_start    ( fm_done) ,
        .load_done    ( fm_done      ) ,
        .ctrl_start   ( load_start[10] ) , // input
        .ctrl_done    ( rd_done[10]      ) , // output
        .ctrl_offset  ( rd_addr[10]      ) , // input [C_ADDR_WIDTH-1:0]
        .ctrl_length  ( rd_length[10]    ) , // input [C_LENGTH_WIDTH-1:0]
        // AXI4 master interface                             
        .arvalid      ( m10_axi_gmem_ARVALID ) , // output
        .arready      ( m10_axi_gmem_ARREADY ) , // input
        .araddr       ( m10_axi_gmem_ARADDR  ) , // output [C_ADDR_WIDTH-1:0]
        .arid         ( m10_axi_gmem_ARID    ) , // output
        .arlen        ( m10_axi_gmem_ARLEN   ) , // output
        .arsize       ( m10_axi_gmem_ARSIZE  ) , // output [2:0]
        .rvalid       ( m10_axi_gmem_RVALID  ) , // input
        .rready       ( m10_axi_gmem_RREADY  ) , // output
        .rdata        ( m10_axi_gmem_RDATA   ) , // input [C_DATA_WIDTH - 1:0]
        .rlast        ( m10_axi_gmem_RLAST   ) , // input
        .rid          ( m10_axi_gmem_RID     ) , // input
        .rresp        ( m10_axi_gmem_RRESP   ) , // input [1:0]
        // FIFO read signals
        .idle         ( rd_channel_idle[10]   ) ,
        .odone        ( rd_done2[10]          ) ,
        .rd_en        ( rd_en[10]             ) , // input
        .rd_data      ( rd_data[10]           ) , // output [C_DATA_WIDTH - 1:0]
        .rd_tvalid_n  ( rd_tvalid_n[10]       ) // output
    );

    krnl_rtl_read_axi #(
    .C_ADDR_WIDTH     ( C_M_AXI_GMEM_ADDR_WIDTH ) ,
    .C_DATA_WIDTH     ( C_M_AXI_GMEM_DATA_WIDTH ) ,
    .C_LENGTH_WIDTH   ( LP_LENGTH_WIDTH         ) ,
    .C_BURST_LEN      ( LP_AXI_BURST_LEN        ) ,
    .C_LOG_BURST_LEN  ( LP_LOG_BURST_LEN        ) ,
    .C_MAX_OUTSTANDING( LP_RD_MAX_OUTSTANDING   )
    )
    axi_read_master_inst11(
        // System signals
        .aclk         ( ap_clk ) , // input
        .areset       ( rd_reset | dev_load_text |  dev_continue | dev_reset ) , // input
        // Control signals 
        .dev_start    ( fm_done) ,
        .load_done    ( fm_done      ) ,
        .ctrl_start   ( load_start[11] ) , // input
        .ctrl_done    ( rd_done[11]      ) , // output
        .ctrl_offset  ( rd_addr[11]      ) , // input [C_ADDR_WIDTH-1:0]
        .ctrl_length  ( rd_length[11]    ) , // input [C_LENGTH_WIDTH-1:0]
        // AXI4 master interface                             
        .arvalid      ( m11_axi_gmem_ARVALID ) , // output
        .arready      ( m11_axi_gmem_ARREADY ) , // input
        .araddr       ( m11_axi_gmem_ARADDR  ) , // output [C_ADDR_WIDTH-1:0]
        .arid         ( m11_axi_gmem_ARID    ) , // output
        .arlen        ( m11_axi_gmem_ARLEN   ) , // output
        .arsize       ( m11_axi_gmem_ARSIZE  ) , // output [2:0]
        .rvalid       ( m11_axi_gmem_RVALID  ) , // input
        .rready       ( m11_axi_gmem_RREADY  ) , // output
        .rdata        ( m11_axi_gmem_RDATA   ) , // input [C_DATA_WIDTH - 1:0]
        .rlast        ( m11_axi_gmem_RLAST   ) , // input
        .rid          ( m11_axi_gmem_RID     ) , // input
        .rresp        ( m11_axi_gmem_RRESP   ) , // input [1:0]
        // FIFO read signals
        .idle         ( rd_channel_idle[11]   ) ,
        .odone        ( rd_done2[11]          ) ,
        .rd_en        ( rd_en[11]             ) , // input
        .rd_data      ( rd_data[11]           ) , // output [C_DATA_WIDTH - 1:0]
        .rd_tvalid_n  ( rd_tvalid_n[11]       ) // output
    );

    krnl_rtl_read_axi #(
    .C_ADDR_WIDTH     ( C_M_AXI_GMEM_ADDR_WIDTH ) ,
    .C_DATA_WIDTH     ( C_M_AXI_GMEM_DATA_WIDTH ) ,
    .C_LENGTH_WIDTH   ( LP_LENGTH_WIDTH         ) ,
    .C_BURST_LEN      ( LP_AXI_BURST_LEN        ) ,
    .C_LOG_BURST_LEN  ( LP_LOG_BURST_LEN        ) ,
    .C_MAX_OUTSTANDING( LP_RD_MAX_OUTSTANDING   )
    )
    axi_read_master_inst12(
        // System signals
        .aclk         ( ap_clk ) , // input
        .areset       ( rd_reset | dev_load_text |  dev_continue | dev_reset ) , // input
        // Control signals 
        .dev_start    ( fm_done) ,
        .load_done    ( fm_done      ) ,
        .ctrl_start   ( load_start[12] ) , // input
        .ctrl_done    ( rd_done[12]      ) , // output
        .ctrl_offset  ( rd_addr[12]      ) , // input [C_ADDR_WIDTH-1:0]
        .ctrl_length  ( rd_length[12]    ) , // input [C_LENGTH_WIDTH-1:0]
        // AXI4 master interface                             
        .arvalid      ( m12_axi_gmem_ARVALID ) , // output
        .arready      ( m12_axi_gmem_ARREADY ) , // input
        .araddr       ( m12_axi_gmem_ARADDR  ) , // output [C_ADDR_WIDTH-1:0]
        .arid         ( m12_axi_gmem_ARID    ) , // output
        .arlen        ( m12_axi_gmem_ARLEN   ) , // output
        .arsize       ( m12_axi_gmem_ARSIZE  ) , // output [2:0]
        .rvalid       ( m12_axi_gmem_RVALID  ) , // input
        .rready       ( m12_axi_gmem_RREADY  ) , // output
        .rdata        ( m12_axi_gmem_RDATA   ) , // input [C_DATA_WIDTH - 1:0]
        .rlast        ( m12_axi_gmem_RLAST   ) , // input
        .rid          ( m12_axi_gmem_RID     ) , // input
        .rresp        ( m12_axi_gmem_RRESP   ) , // input [1:0]
        // FIFO read signals
        .idle         ( rd_channel_idle[12]   ) ,
        .odone        ( rd_done2[12]          ) ,
        .rd_en        ( rd_en[12]             ) , // input
        .rd_data      ( rd_data[12]           ) , // output [C_DATA_WIDTH - 1:0]
        .rd_tvalid_n  ( rd_tvalid_n[12]       ) // output
    );

    krnl_rtl_read_axi #(
    .C_ADDR_WIDTH     ( C_M_AXI_GMEM_ADDR_WIDTH ) ,
    .C_DATA_WIDTH     ( C_M_AXI_GMEM_DATA_WIDTH ) ,
    .C_LENGTH_WIDTH   ( LP_LENGTH_WIDTH         ) ,
    .C_BURST_LEN      ( LP_AXI_BURST_LEN        ) ,
    .C_LOG_BURST_LEN  ( LP_LOG_BURST_LEN        ) ,
    .C_MAX_OUTSTANDING( LP_RD_MAX_OUTSTANDING   )
    )
    axi_read_master_inst13(
        // System signals
        .aclk         ( ap_clk ) , // input
        .areset       ( rd_reset | dev_load_text |  dev_continue | dev_reset ) , // input
        // Control signals 
        .dev_start    ( fm_done) ,
        .load_done    ( fm_done      ) ,
        .ctrl_start   ( load_start[13] ) , // input
        .ctrl_done    ( rd_done[13]      ) , // output
        .ctrl_offset  ( rd_addr[13]      ) , // input [C_ADDR_WIDTH-1:0]
        .ctrl_length  ( rd_length[13]    ) , // input [C_LENGTH_WIDTH-1:0]
        // AXI4 master interface                             
        .arvalid      ( m13_axi_gmem_ARVALID ) , // output
        .arready      ( m13_axi_gmem_ARREADY ) , // input
        .araddr       ( m13_axi_gmem_ARADDR  ) , // output [C_ADDR_WIDTH-1:0]
        .arid         ( m13_axi_gmem_ARID    ) , // output
        .arlen        ( m13_axi_gmem_ARLEN   ) , // output
        .arsize       ( m13_axi_gmem_ARSIZE  ) , // output [2:0]
        .rvalid       ( m13_axi_gmem_RVALID  ) , // input
        .rready       ( m13_axi_gmem_RREADY  ) , // output
        .rdata        ( m13_axi_gmem_RDATA   ) , // input [C_DATA_WIDTH - 1:0]
        .rlast        ( m13_axi_gmem_RLAST   ) , // input
        .rid          ( m13_axi_gmem_RID     ) , // input
        .rresp        ( m13_axi_gmem_RRESP   ) , // input [1:0]
        // FIFO read signals
        .idle         ( rd_channel_idle[13]   ) ,
        .odone        ( rd_done2[13]          ) ,
        .rd_en        ( rd_en[13]             ) , // input
        .rd_data      ( rd_data[13]           ) , // output [C_DATA_WIDTH - 1:0]
        .rd_tvalid_n  ( rd_tvalid_n[13]       ) // output
    );

    krnl_rtl_read_axi #(
    .C_ADDR_WIDTH     ( C_M_AXI_GMEM_ADDR_WIDTH ) ,
    .C_DATA_WIDTH     ( C_M_AXI_GMEM_DATA_WIDTH ) ,
    .C_LENGTH_WIDTH   ( LP_LENGTH_WIDTH         ) ,
    .C_BURST_LEN      ( LP_AXI_BURST_LEN        ) ,
    .C_LOG_BURST_LEN  ( LP_LOG_BURST_LEN        ) ,
    .C_MAX_OUTSTANDING( LP_RD_MAX_OUTSTANDING   )
    )
    axi_read_master_inst14(
        // System signals
        .aclk         ( ap_clk ) , // input
        .areset       ( rd_reset | dev_load_text |  dev_continue | dev_reset ) , // input
        // Control signals 
        .dev_start    ( fm_done) ,
        .load_done    ( fm_done      ) ,
        .ctrl_start   ( load_start[14] ) , // input
        .ctrl_done    ( rd_done[14]      ) , // output
        .ctrl_offset  ( rd_addr[14]      ) , // input [C_ADDR_WIDTH-1:0]
        .ctrl_length  ( rd_length[14]    ) , // input [C_LENGTH_WIDTH-1:0]
        // AXI4 master interface                             
        .arvalid      ( m14_axi_gmem_ARVALID ) , // output
        .arready      ( m14_axi_gmem_ARREADY ) , // input
        .araddr       ( m14_axi_gmem_ARADDR  ) , // output [C_ADDR_WIDTH-1:0]
        .arid         ( m14_axi_gmem_ARID    ) , // output
        .arlen        ( m14_axi_gmem_ARLEN   ) , // output
        .arsize       ( m14_axi_gmem_ARSIZE  ) , // output [2:0]
        .rvalid       ( m14_axi_gmem_RVALID  ) , // input
        .rready       ( m14_axi_gmem_RREADY  ) , // output
        .rdata        ( m14_axi_gmem_RDATA   ) , // input [C_DATA_WIDTH - 1:0]
        .rlast        ( m14_axi_gmem_RLAST   ) , // input
        .rid          ( m14_axi_gmem_RID     ) , // input
        .rresp        ( m14_axi_gmem_RRESP   ) , // input [1:0]
        // FIFO read signals
        .idle         ( rd_channel_idle[14]   ) ,
        .odone        ( rd_done2[14]          ) ,
        .rd_en        ( rd_en[14]             ) , // input
        .rd_data      ( rd_data[14]           ) , // output [C_DATA_WIDTH - 1:0]
        .rd_tvalid_n  ( rd_tvalid_n[14]       ) // output
    );

    krnl_rtl_read_axi #(
    .C_ADDR_WIDTH     ( C_M_AXI_GMEM_ADDR_WIDTH ) ,
    .C_DATA_WIDTH     ( C_M_AXI_GMEM_DATA_WIDTH ) ,
    .C_LENGTH_WIDTH   ( LP_LENGTH_WIDTH         ) ,
    .C_BURST_LEN      ( LP_AXI_BURST_LEN        ) ,
    .C_LOG_BURST_LEN  ( LP_LOG_BURST_LEN        ) ,
    .C_MAX_OUTSTANDING( LP_RD_MAX_OUTSTANDING   )
    )
    axi_read_master_inst15(
        // System signals
        .aclk         ( ap_clk ) , // input
        .areset       ( rd_reset | dev_load_text |  dev_continue | dev_reset ) , // input
        // Control signals 
        .dev_start    ( fm_done) ,
        .load_done    ( fm_done      ) ,
        .ctrl_start   ( load_start[15] ) , // input
        .ctrl_done    ( rd_done[15]      ) , // output
        .ctrl_offset  ( rd_addr[15]      ) , // input [C_ADDR_WIDTH-1:0]
        .ctrl_length  ( rd_length[15]    ) , // input [C_LENGTH_WIDTH-1:0]
        // AXI4 master interface                             
        .arvalid      ( m15_axi_gmem_ARVALID ) , // output
        .arready      ( m15_axi_gmem_ARREADY ) , // input
        .araddr       ( m15_axi_gmem_ARADDR  ) , // output [C_ADDR_WIDTH-1:0]
        .arid         ( m15_axi_gmem_ARID    ) , // output
        .arlen        ( m15_axi_gmem_ARLEN   ) , // output
        .arsize       ( m15_axi_gmem_ARSIZE  ) , // output [2:0]
        .rvalid       ( m15_axi_gmem_RVALID  ) , // input
        .rready       ( m15_axi_gmem_RREADY  ) , // output
        .rdata        ( m15_axi_gmem_RDATA   ) , // input [C_DATA_WIDTH - 1:0]
        .rlast        ( m15_axi_gmem_RLAST   ) , // input
        .rid          ( m15_axi_gmem_RID     ) , // input
        .rresp        ( m15_axi_gmem_RRESP   ) , // input [1:0]
        // FIFO read signals
        .idle         ( rd_channel_idle[15]   ) ,
        .odone        ( rd_done2[15]          ) ,
        .rd_en        ( rd_en[15]             ) , // input
        .rd_data      ( rd_data[15]           ) , // output [C_DATA_WIDTH - 1:0]
        .rd_tvalid_n  ( rd_tvalid_n[15]       ) // output
    );

    krnl_rtl_read_axi #(
    .C_ADDR_WIDTH     ( C_M_AXI_GMEM_ADDR_WIDTH ) ,
    .C_DATA_WIDTH     ( C_M_AXI_GMEM_DATA_WIDTH ) ,
    .C_LENGTH_WIDTH   ( LP_LENGTH_WIDTH         ) ,
    .C_BURST_LEN      ( LP_AXI_BURST_LEN        ) ,
    .C_LOG_BURST_LEN  ( LP_LOG_BURST_LEN        ) ,
    .C_MAX_OUTSTANDING( LP_RD_MAX_OUTSTANDING   )
    )
    axi_read_master_inst16(
        // System signals
        .aclk         ( ap_clk ) , // input
        .areset       ( rd_reset | dev_load_text |  dev_continue | dev_reset ) , // input
        // Control signals 
        .dev_start    ( fm_done) ,
        .load_done    ( fm_done      ) ,
        .ctrl_start   ( load_start[16] ) , // input
        .ctrl_done    ( rd_done[16]      ) , // output
        .ctrl_offset  ( rd_addr[16]      ) , // input [C_ADDR_WIDTH-1:0]
        .ctrl_length  ( rd_length[16]    ) , // input [C_LENGTH_WIDTH-1:0]
        // AXI4 master interface                             
        .arvalid      ( m16_axi_gmem_ARVALID ) , // output
        .arready      ( m16_axi_gmem_ARREADY ) , // input
        .araddr       ( m16_axi_gmem_ARADDR  ) , // output [C_ADDR_WIDTH-1:0]
        .arid         ( m16_axi_gmem_ARID    ) , // output
        .arlen        ( m16_axi_gmem_ARLEN   ) , // output
        .arsize       ( m16_axi_gmem_ARSIZE  ) , // output [2:0]
        .rvalid       ( m16_axi_gmem_RVALID  ) , // input
        .rready       ( m16_axi_gmem_RREADY  ) , // output
        .rdata        ( m16_axi_gmem_RDATA   ) , // input [C_DATA_WIDTH - 1:0]
        .rlast        ( m16_axi_gmem_RLAST   ) , // input
        .rid          ( m16_axi_gmem_RID     ) , // input
        .rresp        ( m16_axi_gmem_RRESP   ) , // input [1:0]
        // FIFO read signals
        .idle         ( rd_channel_idle[16]   ) ,
        .odone        ( rd_done2[16]          ) ,
        .rd_en        ( rd_en[16]             ) , // input
        .rd_data      ( rd_data[16]           ) , // output [C_DATA_WIDTH - 1:0]
        .rd_tvalid_n  ( rd_tvalid_n[16]       ) // output
    );

    krnl_rtl_read_axi #(
    .C_ADDR_WIDTH     ( C_M_AXI_GMEM_ADDR_WIDTH ) ,
    .C_DATA_WIDTH     ( C_M_AXI_GMEM_DATA_WIDTH ) ,
    .C_LENGTH_WIDTH   ( LP_LENGTH_WIDTH         ) ,
    .C_BURST_LEN      ( LP_AXI_BURST_LEN        ) ,
    .C_LOG_BURST_LEN  ( LP_LOG_BURST_LEN        ) ,
    .C_MAX_OUTSTANDING( LP_RD_MAX_OUTSTANDING   )
    )
    axi_read_master_inst17(
        // System signals
        .aclk         ( ap_clk ) , // input
        .areset       ( rd_reset | dev_load_text |  dev_continue | dev_reset ) , // input
        // Control signals 
        .dev_start    ( fm_done) ,
        .load_done    ( fm_done      ) ,
        .ctrl_start   ( load_start[17] ) , // input
        .ctrl_done    ( rd_done[17]      ) , // output
        .ctrl_offset  ( rd_addr[17]      ) , // input [C_ADDR_WIDTH-1:0]
        .ctrl_length  ( rd_length[17]    ) , // input [C_LENGTH_WIDTH-1:0]
        // AXI4 master interface                             
        .arvalid      ( m17_axi_gmem_ARVALID ) , // output
        .arready      ( m17_axi_gmem_ARREADY ) , // input
        .araddr       ( m17_axi_gmem_ARADDR  ) , // output [C_ADDR_WIDTH-1:0]
        .arid         ( m17_axi_gmem_ARID    ) , // output
        .arlen        ( m17_axi_gmem_ARLEN   ) , // output
        .arsize       ( m17_axi_gmem_ARSIZE  ) , // output [2:0]
        .rvalid       ( m17_axi_gmem_RVALID  ) , // input
        .rready       ( m17_axi_gmem_RREADY  ) , // output
        .rdata        ( m17_axi_gmem_RDATA   ) , // input [C_DATA_WIDTH - 1:0]
        .rlast        ( m17_axi_gmem_RLAST   ) , // input
        .rid          ( m17_axi_gmem_RID     ) , // input
        .rresp        ( m17_axi_gmem_RRESP   ) , // input [1:0]
        // FIFO read signals
        .idle         ( rd_channel_idle[17]   ) ,
        .odone        ( rd_done2[17]          ) ,
        .rd_en        ( rd_en[17]             ) , // input
        .rd_data      ( rd_data[17]           ) , // output [C_DATA_WIDTH - 1:0]
        .rd_tvalid_n  ( rd_tvalid_n[17]       ) // output
    );

    krnl_rtl_read_axi #(
    .C_ADDR_WIDTH     ( C_M_AXI_GMEM_ADDR_WIDTH ) ,
    .C_DATA_WIDTH     ( C_M_AXI_GMEM_DATA_WIDTH ) ,
    .C_LENGTH_WIDTH   ( LP_LENGTH_WIDTH         ) ,
    .C_BURST_LEN      ( LP_AXI_BURST_LEN        ) ,
    .C_LOG_BURST_LEN  ( LP_LOG_BURST_LEN        ) ,
    .C_MAX_OUTSTANDING( LP_RD_MAX_OUTSTANDING   )
    )
    axi_read_master_inst18(
        // System signals
        .aclk         ( ap_clk ) , // input
        .areset       ( rd_reset | dev_load_text |  dev_continue | dev_reset ) , // input
        // Control signals 
        .dev_start    ( fm_done) ,
        .load_done    ( fm_done      ) ,
        .ctrl_start   ( load_start[18] ) , // input
        .ctrl_done    ( rd_done[18]      ) , // output
        .ctrl_offset  ( rd_addr[18]      ) , // input [C_ADDR_WIDTH-1:0]
        .ctrl_length  ( rd_length[18]    ) , // input [C_LENGTH_WIDTH-1:0]
        // AXI4 master interface                             
        .arvalid      ( m18_axi_gmem_ARVALID ) , // output
        .arready      ( m18_axi_gmem_ARREADY ) , // input
        .araddr       ( m18_axi_gmem_ARADDR  ) , // output [C_ADDR_WIDTH-1:0]
        .arid         ( m18_axi_gmem_ARID    ) , // output
        .arlen        ( m18_axi_gmem_ARLEN   ) , // output
        .arsize       ( m18_axi_gmem_ARSIZE  ) , // output [2:0]
        .rvalid       ( m18_axi_gmem_RVALID  ) , // input
        .rready       ( m18_axi_gmem_RREADY  ) , // output
        .rdata        ( m18_axi_gmem_RDATA   ) , // input [C_DATA_WIDTH - 1:0]
        .rlast        ( m18_axi_gmem_RLAST   ) , // input
        .rid          ( m18_axi_gmem_RID     ) , // input
        .rresp        ( m18_axi_gmem_RRESP   ) , // input [1:0]
        // FIFO read signals
        .idle         ( rd_channel_idle[18]   ) ,
        .odone        ( rd_done2[18]          ) ,
        .rd_en        ( rd_en[18]             ) , // input
        .rd_data      ( rd_data[18]           ) , // output [C_DATA_WIDTH - 1:0]
        .rd_tvalid_n  ( rd_tvalid_n[18]       ) // output
    );

    krnl_rtl_read_axi #(
    .C_ADDR_WIDTH     ( C_M_AXI_GMEM_ADDR_WIDTH ) ,
    .C_DATA_WIDTH     ( C_M_AXI_GMEM_DATA_WIDTH ) ,
    .C_LENGTH_WIDTH   ( LP_LENGTH_WIDTH         ) ,
    .C_BURST_LEN      ( LP_AXI_BURST_LEN        ) ,
    .C_LOG_BURST_LEN  ( LP_LOG_BURST_LEN        ) ,
    .C_MAX_OUTSTANDING( LP_RD_MAX_OUTSTANDING   )
    )
    axi_read_master_inst19(
        // System signals
        .aclk         ( ap_clk ) , // input
        .areset       ( rd_reset | dev_load_text |  dev_continue | dev_reset ) , // input
        // Control signals 
        .dev_start    ( fm_done) ,
        .load_done    ( fm_done      ) ,
        .ctrl_start   ( load_start[19] ) , // input
        .ctrl_done    ( rd_done[19]      ) , // output
        .ctrl_offset  ( rd_addr[19]      ) , // input [C_ADDR_WIDTH-1:0]
        .ctrl_length  ( rd_length[19]    ) , // input [C_LENGTH_WIDTH-1:0]
        // AXI4 master interface                             
        .arvalid      ( m19_axi_gmem_ARVALID ) , // output
        .arready      ( m19_axi_gmem_ARREADY ) , // input
        .araddr       ( m19_axi_gmem_ARADDR  ) , // output [C_ADDR_WIDTH-1:0]
        .arid         ( m19_axi_gmem_ARID    ) , // output
        .arlen        ( m19_axi_gmem_ARLEN   ) , // output
        .arsize       ( m19_axi_gmem_ARSIZE  ) , // output [2:0]
        .rvalid       ( m19_axi_gmem_RVALID  ) , // input
        .rready       ( m19_axi_gmem_RREADY  ) , // output
        .rdata        ( m19_axi_gmem_RDATA   ) , // input [C_DATA_WIDTH - 1:0]
        .rlast        ( m19_axi_gmem_RLAST   ) , // input
        .rid          ( m19_axi_gmem_RID     ) , // input
        .rresp        ( m19_axi_gmem_RRESP   ) , // input [1:0]
        // FIFO read signals
        .idle         ( rd_channel_idle[19]   ) ,
        .odone        ( rd_done2[19]          ) ,
        .rd_en        ( rd_en[19]             ) , // input
        .rd_data      ( rd_data[19]           ) , // output [C_DATA_WIDTH - 1:0]
        .rd_tvalid_n  ( rd_tvalid_n[19]       ) // output
    );

    krnl_rtl_read_axi #(
    .C_ADDR_WIDTH     ( C_M_AXI_GMEM_ADDR_WIDTH ) ,
    .C_DATA_WIDTH     ( C_M_AXI_GMEM_DATA_WIDTH ) ,
    .C_LENGTH_WIDTH   ( LP_LENGTH_WIDTH         ) ,
    .C_BURST_LEN      ( LP_AXI_BURST_LEN        ) ,
    .C_LOG_BURST_LEN  ( LP_LOG_BURST_LEN        ) ,
    .C_MAX_OUTSTANDING( LP_RD_MAX_OUTSTANDING   )
    )
    axi_read_master_inst20(
        // System signals
        .aclk         ( ap_clk ) , // input
        .areset       ( rd_reset | dev_load_text |  dev_continue | dev_reset ) , // input
        // Control signals 
        .dev_start    ( fm_done) ,
        .load_done    ( fm_done      ) ,
        .ctrl_start   ( load_start[20] ) , // input
        .ctrl_done    ( rd_done[20]      ) , // output
        .ctrl_offset  ( rd_addr[20]      ) , // input [C_ADDR_WIDTH-1:0]
        .ctrl_length  ( rd_length[20]    ) , // input [C_LENGTH_WIDTH-1:0]
        // AXI4 master interface                             
        .arvalid      ( m20_axi_gmem_ARVALID ) , // output
        .arready      ( m20_axi_gmem_ARREADY ) , // input
        .araddr       ( m20_axi_gmem_ARADDR  ) , // output [C_ADDR_WIDTH-1:0]
        .arid         ( m20_axi_gmem_ARID    ) , // output
        .arlen        ( m20_axi_gmem_ARLEN   ) , // output
        .arsize       ( m20_axi_gmem_ARSIZE  ) , // output [2:0]
        .rvalid       ( m20_axi_gmem_RVALID  ) , // input
        .rready       ( m20_axi_gmem_RREADY  ) , // output
        .rdata        ( m20_axi_gmem_RDATA   ) , // input [C_DATA_WIDTH - 1:0]
        .rlast        ( m20_axi_gmem_RLAST   ) , // input
        .rid          ( m20_axi_gmem_RID     ) , // input
        .rresp        ( m20_axi_gmem_RRESP   ) , // input [1:0]
        // FIFO read signals
        .idle         ( rd_channel_idle[20]   ) ,
        .odone        ( rd_done2[20]          ) ,
        .rd_en        ( rd_en[20]             ) , // input
        .rd_data      ( rd_data[20]           ) , // output [C_DATA_WIDTH - 1:0]
        .rd_tvalid_n  ( rd_tvalid_n[20]       ) // output
    );

    krnl_rtl_read_axi #(
    .C_ADDR_WIDTH     ( C_M_AXI_GMEM_ADDR_WIDTH ) ,
    .C_DATA_WIDTH     ( C_M_AXI_GMEM_DATA_WIDTH ) ,
    .C_LENGTH_WIDTH   ( LP_LENGTH_WIDTH         ) ,
    .C_BURST_LEN      ( LP_AXI_BURST_LEN        ) ,
    .C_LOG_BURST_LEN  ( LP_LOG_BURST_LEN        ) ,
    .C_MAX_OUTSTANDING( LP_RD_MAX_OUTSTANDING   )
    )
    axi_read_master_inst21(
        // System signals
        .aclk         ( ap_clk ) , // input
        .areset       ( rd_reset | dev_load_text |  dev_continue | dev_reset ) , // input
        // Control signals 
        .dev_start    ( fm_done) ,
        .load_done    ( fm_done      ) ,
        .ctrl_start   ( load_start[21] ) , // input
        .ctrl_done    ( rd_done[21]      ) , // output
        .ctrl_offset  ( rd_addr[21]      ) , // input [C_ADDR_WIDTH-1:0]
        .ctrl_length  ( rd_length[21]    ) , // input [C_LENGTH_WIDTH-1:0]
        // AXI4 master interface                             
        .arvalid      ( m21_axi_gmem_ARVALID ) , // output
        .arready      ( m21_axi_gmem_ARREADY ) , // input
        .araddr       ( m21_axi_gmem_ARADDR  ) , // output [C_ADDR_WIDTH-1:0]
        .arid         ( m21_axi_gmem_ARID    ) , // output
        .arlen        ( m21_axi_gmem_ARLEN   ) , // output
        .arsize       ( m21_axi_gmem_ARSIZE  ) , // output [2:0]
        .rvalid       ( m21_axi_gmem_RVALID  ) , // input
        .rready       ( m21_axi_gmem_RREADY  ) , // output
        .rdata        ( m21_axi_gmem_RDATA   ) , // input [C_DATA_WIDTH - 1:0]
        .rlast        ( m21_axi_gmem_RLAST   ) , // input
        .rid          ( m21_axi_gmem_RID     ) , // input
        .rresp        ( m21_axi_gmem_RRESP   ) , // input [1:0]
        // FIFO read signals
        .idle         ( rd_channel_idle[21]   ) ,
        .odone        ( rd_done2[21]          ) ,
        .rd_en        ( rd_en[21]             ) , // input
        .rd_data      ( rd_data[21]           ) , // output [C_DATA_WIDTH - 1:0]
        .rd_tvalid_n  ( rd_tvalid_n[21]       ) // output
    );

    krnl_rtl_read_axi #(
    .C_ADDR_WIDTH     ( C_M_AXI_GMEM_ADDR_WIDTH ) ,
    .C_DATA_WIDTH     ( C_M_AXI_GMEM_DATA_WIDTH ) ,
    .C_LENGTH_WIDTH   ( LP_LENGTH_WIDTH         ) ,
    .C_BURST_LEN      ( LP_AXI_BURST_LEN        ) ,
    .C_LOG_BURST_LEN  ( LP_LOG_BURST_LEN        ) ,
    .C_MAX_OUTSTANDING( LP_RD_MAX_OUTSTANDING   )
    )
    axi_read_master_inst22(
        // System signals
        .aclk         ( ap_clk ) , // input
        .areset       ( rd_reset | dev_load_text |  dev_continue | dev_reset ) , // input
        // Control signals 
        .dev_start    ( fm_done) ,
        .load_done    ( fm_done      ) ,
        .ctrl_start   ( load_start[22] ) , // input
        .ctrl_done    ( rd_done[22]      ) , // output
        .ctrl_offset  ( rd_addr[22]      ) , // input [C_ADDR_WIDTH-1:0]
        .ctrl_length  ( rd_length[22]    ) , // input [C_LENGTH_WIDTH-1:0]
        // AXI4 master interface                             
        .arvalid      ( m22_axi_gmem_ARVALID ) , // output
        .arready      ( m22_axi_gmem_ARREADY ) , // input
        .araddr       ( m22_axi_gmem_ARADDR  ) , // output [C_ADDR_WIDTH-1:0]
        .arid         ( m22_axi_gmem_ARID    ) , // output
        .arlen        ( m22_axi_gmem_ARLEN   ) , // output
        .arsize       ( m22_axi_gmem_ARSIZE  ) , // output [2:0]
        .rvalid       ( m22_axi_gmem_RVALID  ) , // input
        .rready       ( m22_axi_gmem_RREADY  ) , // output
        .rdata        ( m22_axi_gmem_RDATA   ) , // input [C_DATA_WIDTH - 1:0]
        .rlast        ( m22_axi_gmem_RLAST   ) , // input
        .rid          ( m22_axi_gmem_RID     ) , // input
        .rresp        ( m22_axi_gmem_RRESP   ) , // input [1:0]
        // FIFO read signals
        .idle         ( rd_channel_idle[22]   ) ,
        .odone        ( rd_done2[22]          ) ,
        .rd_en        ( rd_en[22]             ) , // input
        .rd_data      ( rd_data[22]           ) , // output [C_DATA_WIDTH - 1:0]
        .rd_tvalid_n  ( rd_tvalid_n[22]       ) // output
    );

    krnl_rtl_read_axi #(
    .C_ADDR_WIDTH     ( C_M_AXI_GMEM_ADDR_WIDTH ) ,
    .C_DATA_WIDTH     ( C_M_AXI_GMEM_DATA_WIDTH ) ,
    .C_LENGTH_WIDTH   ( LP_LENGTH_WIDTH         ) ,
    .C_BURST_LEN      ( LP_AXI_BURST_LEN        ) ,
    .C_LOG_BURST_LEN  ( LP_LOG_BURST_LEN        ) ,
    .C_MAX_OUTSTANDING( LP_RD_MAX_OUTSTANDING   )
    )
    axi_read_master_inst23(
        // System signals
        .aclk         ( ap_clk ) , // input
        .areset       ( rd_reset | dev_load_text |  dev_continue | dev_reset ) , // input
        // Control signals 
        .dev_start    ( fm_done) ,
        .load_done    ( fm_done      ) ,
        .ctrl_start   ( load_start[23] ) , // input
        .ctrl_done    ( rd_done[23]      ) , // output
        .ctrl_offset  ( rd_addr[23]      ) , // input [C_ADDR_WIDTH-1:0]
        .ctrl_length  ( rd_length[23]    ) , // input [C_LENGTH_WIDTH-1:0]
        // AXI4 master interface                             
        .arvalid      ( m23_axi_gmem_ARVALID ) , // output
        .arready      ( m23_axi_gmem_ARREADY ) , // input
        .araddr       ( m23_axi_gmem_ARADDR  ) , // output [C_ADDR_WIDTH-1:0]
        .arid         ( m23_axi_gmem_ARID    ) , // output
        .arlen        ( m23_axi_gmem_ARLEN   ) , // output
        .arsize       ( m23_axi_gmem_ARSIZE  ) , // output [2:0]
        .rvalid       ( m23_axi_gmem_RVALID  ) , // input
        .rready       ( m23_axi_gmem_RREADY  ) , // output
        .rdata        ( m23_axi_gmem_RDATA   ) , // input [C_DATA_WIDTH - 1:0]
        .rlast        ( m23_axi_gmem_RLAST   ) , // input
        .rid          ( m23_axi_gmem_RID     ) , // input
        .rresp        ( m23_axi_gmem_RRESP   ) , // input [1:0]
        // FIFO read signals
        .idle         ( rd_channel_idle[23]   ) ,
        .odone        ( rd_done2[23]          ) ,
        .rd_en        ( rd_en[23]             ) , // input
        .rd_data      ( rd_data[23]           ) , // output [C_DATA_WIDTH - 1:0]
        .rd_tvalid_n  ( rd_tvalid_n[23]       ) // output
    );

    krnl_rtl_read_axi #(
    .C_ADDR_WIDTH     ( C_M_AXI_GMEM_ADDR_WIDTH ) ,
    .C_DATA_WIDTH     ( C_M_AXI_GMEM_DATA_WIDTH ) ,
    .C_LENGTH_WIDTH   ( LP_LENGTH_WIDTH         ) ,
    .C_BURST_LEN      ( LP_AXI_BURST_LEN        ) ,
    .C_LOG_BURST_LEN  ( LP_LOG_BURST_LEN        ) ,
    .C_MAX_OUTSTANDING( LP_RD_MAX_OUTSTANDING   )
    )
    axi_read_master_inst24(
        // System signals
        .aclk         ( ap_clk ) , // input
        .areset       ( rd_reset | dev_load_text |  dev_continue | dev_reset ) , // input
        // Control signals 
        .dev_start    ( fm_done) ,
        .load_done    ( fm_done      ) ,
        .ctrl_start   ( load_start[24] ) , // input
        .ctrl_done    ( rd_done[24]      ) , // output
        .ctrl_offset  ( rd_addr[24]      ) , // input [C_ADDR_WIDTH-1:0]
        .ctrl_length  ( rd_length[24]    ) , // input [C_LENGTH_WIDTH-1:0]
        // AXI4 master interface                             
        .arvalid      ( m24_axi_gmem_ARVALID ) , // output
        .arready      ( m24_axi_gmem_ARREADY ) , // input
        .araddr       ( m24_axi_gmem_ARADDR  ) , // output [C_ADDR_WIDTH-1:0]
        .arid         ( m24_axi_gmem_ARID    ) , // output
        .arlen        ( m24_axi_gmem_ARLEN   ) , // output
        .arsize       ( m24_axi_gmem_ARSIZE  ) , // output [2:0]
        .rvalid       ( m24_axi_gmem_RVALID  ) , // input
        .rready       ( m24_axi_gmem_RREADY  ) , // output
        .rdata        ( m24_axi_gmem_RDATA   ) , // input [C_DATA_WIDTH - 1:0]
        .rlast        ( m24_axi_gmem_RLAST   ) , // input
        .rid          ( m24_axi_gmem_RID     ) , // input
        .rresp        ( m24_axi_gmem_RRESP   ) , // input [1:0]
        // FIFO read signals
        .idle         ( rd_channel_idle[24]   ) ,
        .odone        ( rd_done2[24]          ) ,
        .rd_en        ( rd_en[24]             ) , // input
        .rd_data      ( rd_data[24]           ) , // output [C_DATA_WIDTH - 1:0]
        .rd_tvalid_n  ( rd_tvalid_n[24]       ) // output
    );

    krnl_rtl_read_axi #(
    .C_ADDR_WIDTH     ( C_M_AXI_GMEM_ADDR_WIDTH ) ,
    .C_DATA_WIDTH     ( C_M_AXI_GMEM_DATA_WIDTH ) ,
    .C_LENGTH_WIDTH   ( LP_LENGTH_WIDTH         ) ,
    .C_BURST_LEN      ( LP_AXI_BURST_LEN        ) ,
    .C_LOG_BURST_LEN  ( LP_LOG_BURST_LEN        ) ,
    .C_MAX_OUTSTANDING( LP_RD_MAX_OUTSTANDING   )
    )
    axi_read_master_inst25(
        // System signals
        .aclk         ( ap_clk ) , // input
        .areset       ( rd_reset | dev_load_text |  dev_continue | dev_reset ) , // input
        // Control signals 
        .dev_start    ( fm_done) ,
        .load_done    ( fm_done      ) ,
        .ctrl_start   ( load_start[25] ) , // input
        .ctrl_done    ( rd_done[25]      ) , // output
        .ctrl_offset  ( rd_addr[25]      ) , // input [C_ADDR_WIDTH-1:0]
        .ctrl_length  ( rd_length[25]    ) , // input [C_LENGTH_WIDTH-1:0]
        // AXI4 master interface                             
        .arvalid      ( m25_axi_gmem_ARVALID ) , // output
        .arready      ( m25_axi_gmem_ARREADY ) , // input
        .araddr       ( m25_axi_gmem_ARADDR  ) , // output [C_ADDR_WIDTH-1:0]
        .arid         ( m25_axi_gmem_ARID    ) , // output
        .arlen        ( m25_axi_gmem_ARLEN   ) , // output
        .arsize       ( m25_axi_gmem_ARSIZE  ) , // output [2:0]
        .rvalid       ( m25_axi_gmem_RVALID  ) , // input
        .rready       ( m25_axi_gmem_RREADY  ) , // output
        .rdata        ( m25_axi_gmem_RDATA   ) , // input [C_DATA_WIDTH - 1:0]
        .rlast        ( m25_axi_gmem_RLAST   ) , // input
        .rid          ( m25_axi_gmem_RID     ) , // input
        .rresp        ( m25_axi_gmem_RRESP   ) , // input [1:0]
        // FIFO read signals
        .idle         ( rd_channel_idle[25]   ) ,
        .odone        ( rd_done2[25]          ) ,
        .rd_en        ( rd_en[25]             ) , // input
        .rd_data      ( rd_data[25]           ) , // output [C_DATA_WIDTH - 1:0]
        .rd_tvalid_n  ( rd_tvalid_n[25]       ) // output
    );

    krnl_rtl_read_axi #(
    .C_ADDR_WIDTH     ( C_M_AXI_GMEM_ADDR_WIDTH ) ,
    .C_DATA_WIDTH     ( C_M_AXI_GMEM_DATA_WIDTH ) ,
    .C_LENGTH_WIDTH   ( LP_LENGTH_WIDTH         ) ,
    .C_BURST_LEN      ( LP_AXI_BURST_LEN        ) ,
    .C_LOG_BURST_LEN  ( LP_LOG_BURST_LEN        ) ,
    .C_MAX_OUTSTANDING( LP_RD_MAX_OUTSTANDING   )
    )
    axi_read_master_inst26(
        // System signals
        .aclk         ( ap_clk ) , // input
        .areset       ( rd_reset | dev_load_text |  dev_continue | dev_reset ) , // input
        // Control signals 
        .dev_start    ( fm_done) ,
        .load_done    ( fm_done      ) ,
        .ctrl_start   ( load_start[26] ) , // input
        .ctrl_done    ( rd_done[26]      ) , // output
        .ctrl_offset  ( rd_addr[26]      ) , // input [C_ADDR_WIDTH-1:0]
        .ctrl_length  ( rd_length[26]    ) , // input [C_LENGTH_WIDTH-1:0]
        // AXI4 master interface                             
        .arvalid      ( m26_axi_gmem_ARVALID ) , // output
        .arready      ( m26_axi_gmem_ARREADY ) , // input
        .araddr       ( m26_axi_gmem_ARADDR  ) , // output [C_ADDR_WIDTH-1:0]
        .arid         ( m26_axi_gmem_ARID    ) , // output
        .arlen        ( m26_axi_gmem_ARLEN   ) , // output
        .arsize       ( m26_axi_gmem_ARSIZE  ) , // output [2:0]
        .rvalid       ( m26_axi_gmem_RVALID  ) , // input
        .rready       ( m26_axi_gmem_RREADY  ) , // output
        .rdata        ( m26_axi_gmem_RDATA   ) , // input [C_DATA_WIDTH - 1:0]
        .rlast        ( m26_axi_gmem_RLAST   ) , // input
        .rid          ( m26_axi_gmem_RID     ) , // input
        .rresp        ( m26_axi_gmem_RRESP   ) , // input [1:0]
        // FIFO read signals
        .idle         ( rd_channel_idle[26]   ) ,
        .odone        ( rd_done2[26]          ) ,
        .rd_en        ( rd_en[26]             ) , // input
        .rd_data      ( rd_data[26]           ) , // output [C_DATA_WIDTH - 1:0]
        .rd_tvalid_n  ( rd_tvalid_n[26]       ) // output
    );

    krnl_rtl_read_axi #(
    .C_ADDR_WIDTH     ( C_M_AXI_GMEM_ADDR_WIDTH ) ,
    .C_DATA_WIDTH     ( C_M_AXI_GMEM_DATA_WIDTH ) ,
    .C_LENGTH_WIDTH   ( LP_LENGTH_WIDTH         ) ,
    .C_BURST_LEN      ( LP_AXI_BURST_LEN        ) ,
    .C_LOG_BURST_LEN  ( LP_LOG_BURST_LEN        ) ,
    .C_MAX_OUTSTANDING( LP_RD_MAX_OUTSTANDING   )
    )
    axi_read_master_inst27(
        // System signals
        .aclk         ( ap_clk ) , // input
        .areset       ( rd_reset | dev_load_text |  dev_continue | dev_reset ) , // input
        // Control signals 
        .dev_start    ( fm_done) ,
        .load_done    ( fm_done      ) ,
        .ctrl_start   ( load_start[27] ) , // input
        .ctrl_done    ( rd_done[27]      ) , // output
        .ctrl_offset  ( rd_addr[27]      ) , // input [C_ADDR_WIDTH-1:0]
        .ctrl_length  ( rd_length[27]    ) , // input [C_LENGTH_WIDTH-1:0]
        // AXI4 master interface                             
        .arvalid      ( m27_axi_gmem_ARVALID ) , // output
        .arready      ( m27_axi_gmem_ARREADY ) , // input
        .araddr       ( m27_axi_gmem_ARADDR  ) , // output [C_ADDR_WIDTH-1:0]
        .arid         ( m27_axi_gmem_ARID    ) , // output
        .arlen        ( m27_axi_gmem_ARLEN   ) , // output
        .arsize       ( m27_axi_gmem_ARSIZE  ) , // output [2:0]
        .rvalid       ( m27_axi_gmem_RVALID  ) , // input
        .rready       ( m27_axi_gmem_RREADY  ) , // output
        .rdata        ( m27_axi_gmem_RDATA   ) , // input [C_DATA_WIDTH - 1:0]
        .rlast        ( m27_axi_gmem_RLAST   ) , // input
        .rid          ( m27_axi_gmem_RID     ) , // input
        .rresp        ( m27_axi_gmem_RRESP   ) , // input [1:0]
        // FIFO read signals
        .idle         ( rd_channel_idle[27]   ) ,
        .odone        ( rd_done2[27]          ) ,
        .rd_en        ( rd_en[27]             ) , // input
        .rd_data      ( rd_data[27]           ) , // output [C_DATA_WIDTH - 1:0]
        .rd_tvalid_n  ( rd_tvalid_n[27]       ) // output
    );

    krnl_rtl_read_axi #(
    .C_ADDR_WIDTH     ( C_M_AXI_GMEM_ADDR_WIDTH ) ,
    .C_DATA_WIDTH     ( C_M_AXI_GMEM_DATA_WIDTH ) ,
    .C_LENGTH_WIDTH   ( LP_LENGTH_WIDTH         ) ,
    .C_BURST_LEN      ( LP_AXI_BURST_LEN        ) ,
    .C_LOG_BURST_LEN  ( LP_LOG_BURST_LEN        ) ,
    .C_MAX_OUTSTANDING( LP_RD_MAX_OUTSTANDING   )
    )
    axi_read_master_inst28(
        // System signals
        .aclk         ( ap_clk ) , // input
        .areset       ( rd_reset | dev_load_text |  dev_continue | dev_reset ) , // input
        // Control signals 
        .dev_start    ( fm_done) ,
        .load_done    ( fm_done      ) ,
        .ctrl_start   ( load_start[28] ) , // input
        .ctrl_done    ( rd_done[28]      ) , // output
        .ctrl_offset  ( rd_addr[28]      ) , // input [C_ADDR_WIDTH-1:0]
        .ctrl_length  ( rd_length[28]    ) , // input [C_LENGTH_WIDTH-1:0]
        // AXI4 master interface                             
        .arvalid      ( m28_axi_gmem_ARVALID ) , // output
        .arready      ( m28_axi_gmem_ARREADY ) , // input
        .araddr       ( m28_axi_gmem_ARADDR  ) , // output [C_ADDR_WIDTH-1:0]
        .arid         ( m28_axi_gmem_ARID    ) , // output
        .arlen        ( m28_axi_gmem_ARLEN   ) , // output
        .arsize       ( m28_axi_gmem_ARSIZE  ) , // output [2:0]
        .rvalid       ( m28_axi_gmem_RVALID  ) , // input
        .rready       ( m28_axi_gmem_RREADY  ) , // output
        .rdata        ( m28_axi_gmem_RDATA   ) , // input [C_DATA_WIDTH - 1:0]
        .rlast        ( m28_axi_gmem_RLAST   ) , // input
        .rid          ( m28_axi_gmem_RID     ) , // input
        .rresp        ( m28_axi_gmem_RRESP   ) , // input [1:0]
        // FIFO read signals
        .idle         ( rd_channel_idle[28]   ) ,
        .odone        ( rd_done2[28]          ) ,
        .rd_en        ( rd_en[28]             ) , // input
        .rd_data      ( rd_data[28]           ) , // output [C_DATA_WIDTH - 1:0]
        .rd_tvalid_n  ( rd_tvalid_n[28]       ) // output
    );

    krnl_rtl_read_axi #(
    .C_ADDR_WIDTH     ( C_M_AXI_GMEM_ADDR_WIDTH ) ,
    .C_DATA_WIDTH     ( C_M_AXI_GMEM_DATA_WIDTH ) ,
    .C_LENGTH_WIDTH   ( LP_LENGTH_WIDTH         ) ,
    .C_BURST_LEN      ( LP_AXI_BURST_LEN        ) ,
    .C_LOG_BURST_LEN  ( LP_LOG_BURST_LEN        ) ,
    .C_MAX_OUTSTANDING( LP_RD_MAX_OUTSTANDING   )
    )
    axi_read_master_inst29(
        // System signals
        .aclk         ( ap_clk ) , // input
        .areset       ( rd_reset | dev_load_text |  dev_continue | dev_reset ) , // input
        // Control signals 
        .dev_start    ( fm_done) ,
        .load_done    ( fm_done      ) ,
        .ctrl_start   ( load_start[29] ) , // input
        .ctrl_done    ( rd_done[29]      ) , // output
        .ctrl_offset  ( rd_addr[29]      ) , // input [C_ADDR_WIDTH-1:0]
        .ctrl_length  ( rd_length[29]    ) , // input [C_LENGTH_WIDTH-1:0]
        // AXI4 master interface                             
        .arvalid      ( m29_axi_gmem_ARVALID ) , // output
        .arready      ( m29_axi_gmem_ARREADY ) , // input
        .araddr       ( m29_axi_gmem_ARADDR  ) , // output [C_ADDR_WIDTH-1:0]
        .arid         ( m29_axi_gmem_ARID    ) , // output
        .arlen        ( m29_axi_gmem_ARLEN   ) , // output
        .arsize       ( m29_axi_gmem_ARSIZE  ) , // output [2:0]
        .rvalid       ( m29_axi_gmem_RVALID  ) , // input
        .rready       ( m29_axi_gmem_RREADY  ) , // output
        .rdata        ( m29_axi_gmem_RDATA   ) , // input [C_DATA_WIDTH - 1:0]
        .rlast        ( m29_axi_gmem_RLAST   ) , // input
        .rid          ( m29_axi_gmem_RID     ) , // input
        .rresp        ( m29_axi_gmem_RRESP   ) , // input [1:0]
        // FIFO read signals
        .idle         ( rd_channel_idle[29]   ) ,
        .odone        ( rd_done2[29]          ) ,
        .rd_en        ( rd_en[29]             ) , // input
        .rd_data      ( rd_data[29]           ) , // output [C_DATA_WIDTH - 1:0]
        .rd_tvalid_n  ( rd_tvalid_n[29]       ) // output
    );

    krnl_rtl_read_axi #(
    .C_ADDR_WIDTH     ( C_M_AXI_GMEM_ADDR_WIDTH ) ,
    .C_DATA_WIDTH     ( C_M_AXI_GMEM_DATA_WIDTH ) ,
    .C_LENGTH_WIDTH   ( LP_LENGTH_WIDTH         ) ,
    .C_BURST_LEN      ( LP_AXI_BURST_LEN        ) ,
    .C_LOG_BURST_LEN  ( LP_LOG_BURST_LEN        ) ,
    .C_MAX_OUTSTANDING( LP_RD_MAX_OUTSTANDING   )
    )
    axi_read_master_inst30(
        // System signals
        .aclk         ( ap_clk ) , // input
        .areset       ( rd_reset | dev_load_text |  dev_continue | dev_reset ) , // input
        // Control signals 
        .dev_start    ( fm_done) ,
        .load_done    ( fm_done      ) ,
        .ctrl_start   ( load_start[30] ) , // input
        .ctrl_done    ( rd_done[30]      ) , // output
        .ctrl_offset  ( rd_addr[30]      ) , // input [C_ADDR_WIDTH-1:0]
        .ctrl_length  ( rd_length[30]    ) , // input [C_LENGTH_WIDTH-1:0]
        // AXI4 master interface                             
        .arvalid      ( m30_axi_gmem_ARVALID ) , // output
        .arready      ( m30_axi_gmem_ARREADY ) , // input
        .araddr       ( m30_axi_gmem_ARADDR  ) , // output [C_ADDR_WIDTH-1:0]
        .arid         ( m30_axi_gmem_ARID    ) , // output
        .arlen        ( m30_axi_gmem_ARLEN   ) , // output
        .arsize       ( m30_axi_gmem_ARSIZE  ) , // output [2:0]
        .rvalid       ( m30_axi_gmem_RVALID  ) , // input
        .rready       ( m30_axi_gmem_RREADY  ) , // output
        .rdata        ( m30_axi_gmem_RDATA   ) , // input [C_DATA_WIDTH - 1:0]
        .rlast        ( m30_axi_gmem_RLAST   ) , // input
        .rid          ( m30_axi_gmem_RID     ) , // input
        .rresp        ( m30_axi_gmem_RRESP   ) , // input [1:0]
        // FIFO read signals
        .idle         ( rd_channel_idle[30]   ) ,
        .odone        ( rd_done2[30]          ) ,
        .rd_en        ( rd_en[30]             ) , // input
        .rd_data      ( rd_data[30]           ) , // output [C_DATA_WIDTH - 1:0]
        .rd_tvalid_n  ( rd_tvalid_n[30]       ) // output
    );

    krnl_rtl_read_axi #(
    .C_ADDR_WIDTH     ( C_M_AXI_GMEM_ADDR_WIDTH ) ,
    .C_DATA_WIDTH     ( C_M_AXI_GMEM_DATA_WIDTH ) ,
    .C_LENGTH_WIDTH   ( LP_LENGTH_WIDTH         ) ,
    .C_BURST_LEN      ( LP_AXI_BURST_LEN        ) ,
    .C_LOG_BURST_LEN  ( LP_LOG_BURST_LEN        ) ,
    .C_MAX_OUTSTANDING( LP_RD_MAX_OUTSTANDING   )
    )
    axi_read_master_inst31(
        // System signals
        .aclk         ( ap_clk ) , // input
        .areset       ( rd_reset | dev_load_text |  dev_continue | dev_reset ) , // input
        // Control signals 
        .dev_start    ( fm_done) ,
        .load_done    ( fm_done      ) ,
        .ctrl_start   ( load_start[31] ) , // input
        .ctrl_done    ( rd_done[31]      ) , // output
        .ctrl_offset  ( rd_addr[31]      ) , // input [C_ADDR_WIDTH-1:0]
        .ctrl_length  ( rd_length[31]    ) , // input [C_LENGTH_WIDTH-1:0]
        // AXI4 master interface                             
        .arvalid      ( m31_axi_gmem_ARVALID ) , // output
        .arready      ( m31_axi_gmem_ARREADY ) , // input
        .araddr       ( m31_axi_gmem_ARADDR  ) , // output [C_ADDR_WIDTH-1:0]
        .arid         ( m31_axi_gmem_ARID    ) , // output
        .arlen        ( m31_axi_gmem_ARLEN   ) , // output
        .arsize       ( m31_axi_gmem_ARSIZE  ) , // output [2:0]
        .rvalid       ( m31_axi_gmem_RVALID  ) , // input
        .rready       ( m31_axi_gmem_RREADY  ) , // output
        .rdata        ( m31_axi_gmem_RDATA   ) , // input [C_DATA_WIDTH - 1:0]
        .rlast        ( m31_axi_gmem_RLAST   ) , // input
        .rid          ( m31_axi_gmem_RID     ) , // input
        .rresp        ( m31_axi_gmem_RRESP   ) , // input [1:0]
        // FIFO read signals
        .idle         ( rd_channel_idle[31]   ) ,
        .odone        ( rd_done2[31]          ) ,
        .rd_en        ( rd_en[31]             ) , // input
        .rd_data      ( rd_data[31]           ) , // output [C_DATA_WIDTH - 1:0]
        .rd_tvalid_n  ( rd_tvalid_n[31]       ) // output
    );

    tsp_top tsp_core(
        .ICLK           ( ap_clk             ) ,
        .IRESET         ( areset | dev_reset |  dev_continue) ,
        .ICONTINUE      ( dev_continue       ) ,
        .IRESETTEXT     ( dev_load_text      ) ,
        .IOVERLAP       ( fm_overlap         ) ,
        // 32 channels 64-bits (update text)
        .ITEXT0_DATA    ( rd_data[0] ) ,
        .ITEXT1_DATA    ( rd_data[1] ) ,
        .ITEXT2_DATA    ( rd_data[2] ) ,
        .ITEXT3_DATA    ( rd_data[3] ) ,
        .ITEXT4_DATA    ( rd_data[4] ) ,
        .ITEXT5_DATA    ( rd_data[5] ) ,
        .ITEXT6_DATA    ( rd_data[6] ) ,
        .ITEXT7_DATA    ( rd_data[7] ) ,
        .ITEXT8_DATA    ( rd_data[8] ) ,
        .ITEXT9_DATA    ( rd_data[9] ) ,
        .ITEXT10_DATA   ( rd_data[10] ) ,
        .ITEXT11_DATA   ( rd_data[11] ) ,
        .ITEXT12_DATA   ( rd_data[12] ) ,
        .ITEXT13_DATA   ( rd_data[13] ) ,
        .ITEXT14_DATA   ( rd_data[14] ) ,
        .ITEXT15_DATA   ( rd_data[15] ) ,
        .ITEXT16_DATA   ( rd_data[16] ) ,
        .ITEXT17_DATA   ( rd_data[17] ) ,
        .ITEXT18_DATA   ( rd_data[18] ) ,
        .ITEXT19_DATA   ( rd_data[19] ) ,
        .ITEXT20_DATA   ( rd_data[20] ) ,
        .ITEXT21_DATA   ( rd_data[21] ) ,
        .ITEXT22_DATA   ( rd_data[22] ) ,
        .ITEXT23_DATA   ( rd_data[23] ) ,
        .ITEXT24_DATA   ( rd_data[24] ) ,
        .ITEXT25_DATA   ( rd_data[25] ) ,
        .ITEXT26_DATA   ( rd_data[26] ) ,
        .ITEXT27_DATA   ( rd_data[27] ) ,
        .ITEXT28_DATA   ( rd_data[28] ) ,
        .ITEXT29_DATA   ( rd_data[29] ) ,
        .ITEXT30_DATA   ( rd_data[30] ) ,
        .ITEXT31_DATA   ( rd_data[31] ) ,
        .ITEXT_WE       ( rd_datavld  ) ,
        .BITSTREAM_RDEN ( bitstream_rden     ) ,
        // Read result port
        .IRDEN              ( result_rden        ) ,
        .ODATA              ( result_data        ) ,
        .ODATAVALID         ( result_valid       ) ,
        .OFULL              (  ) ,
        .OEMPTY             (  ) ,
        .MATCH_COUNT        ( match_count        ) ,
        .MATCH_COUNT_VALID  ( match_count_vld    ) ,
        .BITSTREAM          ( bitstream          ) ,
        .BASH_CODE          (  ) ,
        // Buffer control singnals
        .BUFFER_START       ( dev_start     ) ,
        .BUFFER_BYTEMODE    ( dev_bytemode  ) ,
        .BUFFER_IKEY        ( ikey[13:0]    ) ,
        .BUFFER_WREN        ( ikey_wren     ) ,
        .KEY_LAST           ( key_last      )
    );

    
    assign rd_datavld = ~rd_tvalid_n;
    assign rd_en = rd_datavld;
    
    assign ap_done = key_last;
    assign dev_done = key_last;
    
    assign m00_axi_gmem_AWVALID = 1'b0;
    assign m00_axi_gmem_AWADDR = 64'd0;
    assign m00_axi_gmem_AWLEN  = 8'd0;
    assign m00_axi_gmem_AWSIZE = 3'd0;
    assign m00_axi_gmem_WVALID = 1'b0;
    assign m00_axi_gmem_WDATA = 64'd0;
    assign m00_axi_gmem_WSTRB = 8'd0;
    assign m00_axi_gmem_WLAST = 1'b0;
    assign m00_axi_gmem_BREADY = 1'b0;

    assign m01_axi_gmem_AWVALID = 1'b0;
    assign m01_axi_gmem_AWADDR = 64'd0;
    assign m01_axi_gmem_AWLEN  = 8'd0;
    assign m01_axi_gmem_AWSIZE = 3'd0;
    assign m01_axi_gmem_WVALID = 1'b0;
    assign m01_axi_gmem_WDATA = 64'd0;
    assign m01_axi_gmem_WSTRB = 8'd0;
    assign m01_axi_gmem_WLAST = 1'b0;
    assign m01_axi_gmem_BREADY = 1'b0;

    assign m02_axi_gmem_AWVALID = 1'b0;
    assign m02_axi_gmem_AWADDR = 64'd0;
    assign m02_axi_gmem_AWLEN  = 8'd0;
    assign m02_axi_gmem_AWSIZE = 3'd0;
    assign m02_axi_gmem_WVALID = 1'b0;
    assign m02_axi_gmem_WDATA = 64'd0;
    assign m02_axi_gmem_WSTRB = 8'd0;
    assign m02_axi_gmem_WLAST = 1'b0;
    assign m02_axi_gmem_BREADY = 1'b0;

    assign m03_axi_gmem_AWVALID = 1'b0;
    assign m03_axi_gmem_AWADDR = 64'd0;
    assign m03_axi_gmem_AWLEN  = 8'd0;
    assign m03_axi_gmem_AWSIZE = 3'd0;
    assign m03_axi_gmem_WVALID = 1'b0;
    assign m03_axi_gmem_WDATA = 64'd0;
    assign m03_axi_gmem_WSTRB = 8'd0;
    assign m03_axi_gmem_WLAST = 1'b0;
    assign m03_axi_gmem_BREADY = 1'b0;

    assign m04_axi_gmem_AWVALID = 1'b0;
    assign m04_axi_gmem_AWADDR = 64'd0;
    assign m04_axi_gmem_AWLEN  = 8'd0;
    assign m04_axi_gmem_AWSIZE = 3'd0;
    assign m04_axi_gmem_WVALID = 1'b0;
    assign m04_axi_gmem_WDATA = 64'd0;
    assign m04_axi_gmem_WSTRB = 8'd0;
    assign m04_axi_gmem_WLAST = 1'b0;
    assign m04_axi_gmem_BREADY = 1'b0;

    assign m05_axi_gmem_AWVALID = 1'b0;
    assign m05_axi_gmem_AWADDR = 64'd0;
    assign m05_axi_gmem_AWLEN  = 8'd0;
    assign m05_axi_gmem_AWSIZE = 3'd0;
    assign m05_axi_gmem_WVALID = 1'b0;
    assign m05_axi_gmem_WDATA = 64'd0;
    assign m05_axi_gmem_WSTRB = 8'd0;
    assign m05_axi_gmem_WLAST = 1'b0;
    assign m05_axi_gmem_BREADY = 1'b0;

    assign m06_axi_gmem_AWVALID = 1'b0;
    assign m06_axi_gmem_AWADDR = 64'd0;
    assign m06_axi_gmem_AWLEN  = 8'd0;
    assign m06_axi_gmem_AWSIZE = 3'd0;
    assign m06_axi_gmem_WVALID = 1'b0;
    assign m06_axi_gmem_WDATA = 64'd0;
    assign m06_axi_gmem_WSTRB = 8'd0;
    assign m06_axi_gmem_WLAST = 1'b0;
    assign m06_axi_gmem_BREADY = 1'b0;

    assign m07_axi_gmem_AWVALID = 1'b0;
    assign m07_axi_gmem_AWADDR = 64'd0;
    assign m07_axi_gmem_AWLEN  = 8'd0;
    assign m07_axi_gmem_AWSIZE = 3'd0;
    assign m07_axi_gmem_WVALID = 1'b0;
    assign m07_axi_gmem_WDATA = 64'd0;
    assign m07_axi_gmem_WSTRB = 8'd0;
    assign m07_axi_gmem_WLAST = 1'b0;
    assign m07_axi_gmem_BREADY = 1'b0;

    assign m08_axi_gmem_AWVALID = 1'b0;
    assign m08_axi_gmem_AWADDR = 64'd0;
    assign m08_axi_gmem_AWLEN  = 8'd0;
    assign m08_axi_gmem_AWSIZE = 3'd0;
    assign m08_axi_gmem_WVALID = 1'b0;
    assign m08_axi_gmem_WDATA = 64'd0;
    assign m08_axi_gmem_WSTRB = 8'd0;
    assign m08_axi_gmem_WLAST = 1'b0;
    assign m08_axi_gmem_BREADY = 1'b0;

    assign m09_axi_gmem_AWVALID = 1'b0;
    assign m09_axi_gmem_AWADDR = 64'd0;
    assign m09_axi_gmem_AWLEN  = 8'd0;
    assign m09_axi_gmem_AWSIZE = 3'd0;
    assign m09_axi_gmem_WVALID = 1'b0;
    assign m09_axi_gmem_WDATA = 64'd0;
    assign m09_axi_gmem_WSTRB = 8'd0;
    assign m09_axi_gmem_WLAST = 1'b0;
    assign m09_axi_gmem_BREADY = 1'b0;

    assign m10_axi_gmem_AWVALID = 1'b0;
    assign m10_axi_gmem_AWADDR = 64'd0;
    assign m10_axi_gmem_AWLEN  = 8'd0;
    assign m10_axi_gmem_AWSIZE = 3'd0;
    assign m10_axi_gmem_WVALID = 1'b0;
    assign m10_axi_gmem_WDATA = 64'd0;
    assign m10_axi_gmem_WSTRB = 8'd0;
    assign m10_axi_gmem_WLAST = 1'b0;
    assign m10_axi_gmem_BREADY = 1'b0;

    assign m11_axi_gmem_AWVALID = 1'b0;
    assign m11_axi_gmem_AWADDR = 64'd0;
    assign m11_axi_gmem_AWLEN  = 8'd0;
    assign m11_axi_gmem_AWSIZE = 3'd0;
    assign m11_axi_gmem_WVALID = 1'b0;
    assign m11_axi_gmem_WDATA = 64'd0;
    assign m11_axi_gmem_WSTRB = 8'd0;
    assign m11_axi_gmem_WLAST = 1'b0;
    assign m11_axi_gmem_BREADY = 1'b0;

    assign m12_axi_gmem_AWVALID = 1'b0;
    assign m12_axi_gmem_AWADDR = 64'd0;
    assign m12_axi_gmem_AWLEN  = 8'd0;
    assign m12_axi_gmem_AWSIZE = 3'd0;
    assign m12_axi_gmem_WVALID = 1'b0;
    assign m12_axi_gmem_WDATA = 64'd0;
    assign m12_axi_gmem_WSTRB = 8'd0;
    assign m12_axi_gmem_WLAST = 1'b0;
    assign m12_axi_gmem_BREADY = 1'b0;

    assign m13_axi_gmem_AWVALID = 1'b0;
    assign m13_axi_gmem_AWADDR = 64'd0;
    assign m13_axi_gmem_AWLEN  = 8'd0;
    assign m13_axi_gmem_AWSIZE = 3'd0;
    assign m13_axi_gmem_WVALID = 1'b0;
    assign m13_axi_gmem_WDATA = 64'd0;
    assign m13_axi_gmem_WSTRB = 8'd0;
    assign m13_axi_gmem_WLAST = 1'b0;
    assign m13_axi_gmem_BREADY = 1'b0;

    assign m14_axi_gmem_AWVALID = 1'b0;
    assign m14_axi_gmem_AWADDR = 64'd0;
    assign m14_axi_gmem_AWLEN  = 8'd0;
    assign m14_axi_gmem_AWSIZE = 3'd0;
    assign m14_axi_gmem_WVALID = 1'b0;
    assign m14_axi_gmem_WDATA = 64'd0;
    assign m14_axi_gmem_WSTRB = 8'd0;
    assign m14_axi_gmem_WLAST = 1'b0;
    assign m14_axi_gmem_BREADY = 1'b0;

    assign m15_axi_gmem_AWVALID = 1'b0;
    assign m15_axi_gmem_AWADDR = 64'd0;
    assign m15_axi_gmem_AWLEN  = 8'd0;
    assign m15_axi_gmem_AWSIZE = 3'd0;
    assign m15_axi_gmem_WVALID = 1'b0;
    assign m15_axi_gmem_WDATA = 64'd0;
    assign m15_axi_gmem_WSTRB = 8'd0;
    assign m15_axi_gmem_WLAST = 1'b0;
    assign m15_axi_gmem_BREADY = 1'b0;

    assign m16_axi_gmem_AWVALID = 1'b0;
    assign m16_axi_gmem_AWADDR = 64'd0;
    assign m16_axi_gmem_AWLEN  = 8'd0;
    assign m16_axi_gmem_AWSIZE = 3'd0;
    assign m16_axi_gmem_WVALID = 1'b0;
    assign m16_axi_gmem_WDATA = 64'd0;
    assign m16_axi_gmem_WSTRB = 8'd0;
    assign m16_axi_gmem_WLAST = 1'b0;
    assign m16_axi_gmem_BREADY = 1'b0;

    assign m17_axi_gmem_AWVALID = 1'b0;
    assign m17_axi_gmem_AWADDR = 64'd0;
    assign m17_axi_gmem_AWLEN  = 8'd0;
    assign m17_axi_gmem_AWSIZE = 3'd0;
    assign m17_axi_gmem_WVALID = 1'b0;
    assign m17_axi_gmem_WDATA = 64'd0;
    assign m17_axi_gmem_WSTRB = 8'd0;
    assign m17_axi_gmem_WLAST = 1'b0;
    assign m17_axi_gmem_BREADY = 1'b0;

    assign m18_axi_gmem_AWVALID = 1'b0;
    assign m18_axi_gmem_AWADDR = 64'd0;
    assign m18_axi_gmem_AWLEN  = 8'd0;
    assign m18_axi_gmem_AWSIZE = 3'd0;
    assign m18_axi_gmem_WVALID = 1'b0;
    assign m18_axi_gmem_WDATA = 64'd0;
    assign m18_axi_gmem_WSTRB = 8'd0;
    assign m18_axi_gmem_WLAST = 1'b0;
    assign m18_axi_gmem_BREADY = 1'b0;

    assign m19_axi_gmem_AWVALID = 1'b0;
    assign m19_axi_gmem_AWADDR = 64'd0;
    assign m19_axi_gmem_AWLEN  = 8'd0;
    assign m19_axi_gmem_AWSIZE = 3'd0;
    assign m19_axi_gmem_WVALID = 1'b0;
    assign m19_axi_gmem_WDATA = 64'd0;
    assign m19_axi_gmem_WSTRB = 8'd0;
    assign m19_axi_gmem_WLAST = 1'b0;
    assign m19_axi_gmem_BREADY = 1'b0;

    assign m20_axi_gmem_AWVALID = 1'b0;
    assign m20_axi_gmem_AWADDR = 64'd0;
    assign m20_axi_gmem_AWLEN  = 8'd0;
    assign m20_axi_gmem_AWSIZE = 3'd0;
    assign m20_axi_gmem_WVALID = 1'b0;
    assign m20_axi_gmem_WDATA = 64'd0;
    assign m20_axi_gmem_WSTRB = 8'd0;
    assign m20_axi_gmem_WLAST = 1'b0;
    assign m20_axi_gmem_BREADY = 1'b0;

    assign m21_axi_gmem_AWVALID = 1'b0;
    assign m21_axi_gmem_AWADDR = 64'd0;
    assign m21_axi_gmem_AWLEN  = 8'd0;
    assign m21_axi_gmem_AWSIZE = 3'd0;
    assign m21_axi_gmem_WVALID = 1'b0;
    assign m21_axi_gmem_WDATA = 64'd0;
    assign m21_axi_gmem_WSTRB = 8'd0;
    assign m21_axi_gmem_WLAST = 1'b0;
    assign m21_axi_gmem_BREADY = 1'b0;

    assign m22_axi_gmem_AWVALID = 1'b0;
    assign m22_axi_gmem_AWADDR = 64'd0;
    assign m22_axi_gmem_AWLEN  = 8'd0;
    assign m22_axi_gmem_AWSIZE = 3'd0;
    assign m22_axi_gmem_WVALID = 1'b0;
    assign m22_axi_gmem_WDATA = 64'd0;
    assign m22_axi_gmem_WSTRB = 8'd0;
    assign m22_axi_gmem_WLAST = 1'b0;
    assign m22_axi_gmem_BREADY = 1'b0;

    assign m23_axi_gmem_AWVALID = 1'b0;
    assign m23_axi_gmem_AWADDR = 64'd0;
    assign m23_axi_gmem_AWLEN  = 8'd0;
    assign m23_axi_gmem_AWSIZE = 3'd0;
    assign m23_axi_gmem_WVALID = 1'b0;
    assign m23_axi_gmem_WDATA = 64'd0;
    assign m23_axi_gmem_WSTRB = 8'd0;
    assign m23_axi_gmem_WLAST = 1'b0;
    assign m23_axi_gmem_BREADY = 1'b0;

    assign m24_axi_gmem_AWVALID = 1'b0;
    assign m24_axi_gmem_AWADDR = 64'd0;
    assign m24_axi_gmem_AWLEN  = 8'd0;
    assign m24_axi_gmem_AWSIZE = 3'd0;
    assign m24_axi_gmem_WVALID = 1'b0;
    assign m24_axi_gmem_WDATA = 64'd0;
    assign m24_axi_gmem_WSTRB = 8'd0;
    assign m24_axi_gmem_WLAST = 1'b0;
    assign m24_axi_gmem_BREADY = 1'b0;

    assign m25_axi_gmem_AWVALID = 1'b0;
    assign m25_axi_gmem_AWADDR = 64'd0;
    assign m25_axi_gmem_AWLEN  = 8'd0;
    assign m25_axi_gmem_AWSIZE = 3'd0;
    assign m25_axi_gmem_WVALID = 1'b0;
    assign m25_axi_gmem_WDATA = 64'd0;
    assign m25_axi_gmem_WSTRB = 8'd0;
    assign m25_axi_gmem_WLAST = 1'b0;
    assign m25_axi_gmem_BREADY = 1'b0;

    assign m26_axi_gmem_AWVALID = 1'b0;
    assign m26_axi_gmem_AWADDR = 64'd0;
    assign m26_axi_gmem_AWLEN  = 8'd0;
    assign m26_axi_gmem_AWSIZE = 3'd0;
    assign m26_axi_gmem_WVALID = 1'b0;
    assign m26_axi_gmem_WDATA = 64'd0;
    assign m26_axi_gmem_WSTRB = 8'd0;
    assign m26_axi_gmem_WLAST = 1'b0;
    assign m26_axi_gmem_BREADY = 1'b0;

    assign m27_axi_gmem_AWVALID = 1'b0;
    assign m27_axi_gmem_AWADDR = 64'd0;
    assign m27_axi_gmem_AWLEN  = 8'd0;
    assign m27_axi_gmem_AWSIZE = 3'd0;
    assign m27_axi_gmem_WVALID = 1'b0;
    assign m27_axi_gmem_WDATA = 64'd0;
    assign m27_axi_gmem_WSTRB = 8'd0;
    assign m27_axi_gmem_WLAST = 1'b0;
    assign m27_axi_gmem_BREADY = 1'b0;

    assign m28_axi_gmem_AWVALID = 1'b0;
    assign m28_axi_gmem_AWADDR = 64'd0;
    assign m28_axi_gmem_AWLEN  = 8'd0;
    assign m28_axi_gmem_AWSIZE = 3'd0;
    assign m28_axi_gmem_WVALID = 1'b0;
    assign m28_axi_gmem_WDATA = 64'd0;
    assign m28_axi_gmem_WSTRB = 8'd0;
    assign m28_axi_gmem_WLAST = 1'b0;
    assign m28_axi_gmem_BREADY = 1'b0;

    assign m29_axi_gmem_AWVALID = 1'b0;
    assign m29_axi_gmem_AWADDR = 64'd0;
    assign m29_axi_gmem_AWLEN  = 8'd0;
    assign m29_axi_gmem_AWSIZE = 3'd0;
    assign m29_axi_gmem_WVALID = 1'b0;
    assign m29_axi_gmem_WDATA = 64'd0;
    assign m29_axi_gmem_WSTRB = 8'd0;
    assign m29_axi_gmem_WLAST = 1'b0;
    assign m29_axi_gmem_BREADY = 1'b0;

    assign m30_axi_gmem_AWVALID = 1'b0;
    assign m30_axi_gmem_AWADDR = 64'd0;
    assign m30_axi_gmem_AWLEN  = 8'd0;
    assign m30_axi_gmem_AWSIZE = 3'd0;
    assign m30_axi_gmem_WVALID = 1'b0;
    assign m30_axi_gmem_WDATA = 64'd0;
    assign m30_axi_gmem_WSTRB = 8'd0;
    assign m30_axi_gmem_WLAST = 1'b0;
    assign m30_axi_gmem_BREADY = 1'b0;

    assign m31_axi_gmem_AWVALID = 1'b0;
    assign m31_axi_gmem_AWADDR = 64'd0;
    assign m31_axi_gmem_AWLEN  = 8'd0;
    assign m31_axi_gmem_AWSIZE = 3'd0;
    assign m31_axi_gmem_WVALID = 1'b0;
    assign m31_axi_gmem_WDATA = 64'd0;
    assign m31_axi_gmem_WSTRB = 8'd0;
    assign m31_axi_gmem_WLAST = 1'b0;
    assign m31_axi_gmem_BREADY = 1'b0;

endmodule
